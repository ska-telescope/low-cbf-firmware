----------------------------------------------------------------------------------
-- Company: CSIRO CASS 
-- Engineer: David Humphrey
-- 
-- Create Date: 14.11.2018 11:27:29
-- Module Name: correlatorFBTop25 - Behavioral
-- Description: 
--  Filterbank with 12 FIR taps, 4096 point FFT, critically sampled.
--  Processes 4 parallel signals, each with 8 bit complex data (8 bit real + 8 bit imaginary).
--  This version (with the "25" suffix) refers to the use of 25 bits of precision in the FFT
--  high precision is used to ensure very low bias in the filterbank output (needed to meet the low.CBF 1000 hour noise test).
--  
-- Supporting Code:
--  The Matlab model should be in the directory ../matlab_model
--  Key files:
--   * ../matlab_model/run_correlatorFB.m 
--       Generate input files for the simulation, run the matlab model and compares with simulation output
--   * ../matlab_model/get_rom_coefficients.m
--       Generates ROM data used in the firmware. ROMs are initialised using .coe files.
--       "filtertaps_X.coe" : X runs from 1 to 12, contents of the 12 ROMS used to store the FIR filter taps.
--
--  There is a top level module that can be used to build this in a standalone version 
--   "correlatorFBtesttop.vhd"
-- Structure:
--
--  File Structure
--  --------------
--  Outline of the structure shown below. Excludes .xci files for DSPs, RAMs and ROMs.
--
--    correlatorFBTop.vhd : This file, 4 complex inputs, 12 FIR filter taps, 4096 point FFT.
--        |
--        +-- correlatorFBMem.vhd         : Input memory for the filterbank, 12 blocks of memory chained together. Also holds memory for the coefficients.
--        +-- fb_DSP25.vhd                : 12 TAP FIR filter
--        +-- correlatorFFT25wrapper.vhd  : 4096 point FFT
--                |
--                +-- fft4096_25bit.xci : standard Xilinx 4096 point FFT (4 used).
--
--  TestBench
--  ---------
--  correlatorFB_tb.vhd reads the input data generated by the Matlab model and generates output files for checking by the matlab code.
--
--  Resource Use
--  ------------
--  Approximate resource usage is 
--   LUTs        = 15,607
--   DSPs        = 176
--   Registers   = 27,187
--   BRAMs (36K) = 58
--   URAMs       = 15
--  Note this is about 50% more LUTS and registers as compared with the version that uses 16 bit precision for the FFT (but the same number of DSPs).
-- 
--  Power estimate (Guess based on related measurement on zcu111 board)
--   about 1 W static, 3.5 W dynamic.
--
--  -----------------------------------------------------------------------------------------------
--  Description
--  -----------
--
-- 1. Filterbank Memory
--   The filterbank memory consists of 11 blocks of memory chained together.
--   The read and write addresses are staggered by one clock for each memory, implemented as a 12 sample delay line on
--   the address. This makes the timing easy to meet for the  memory address signals (which would otherwise be high-fanout signals)
--   and also enables use of the adders in the DSPs for the FIR filter.  
--
-- 2. FIR filter
--   The FIR filter uses 12 DSPs for each of the 8 simultaneous samples (4 channels * 2 [real+imaginary]) that are read from the memory.
--   So the FIR filter uses (12 DSPS) * (8 simultaneous samples) = 96 DSPs.
--   The filter is implemented entirely in DSPs. The PCOUT port on the DSP is used to send the result of the multiplication
--   to the next DSP in the chain, where it is added using the adder in the DSP. This scheme requires that the inputs to the
--   12 DSPs are staggered to account for the pipeline stage on the PCOUT port. The staggering is done by controlling the address
--   to the memories as described above.
--
-- 3. 4096 point FFT
--   Standard Xilinx FFT. Some messy logic at the front to account for the delay inserted by the "real-time" mode.
--
-- 4. Reorder memory
--   Data out of the FFT is in bit reversed order. It is stored in a double buffer in order from low to high frequencies,
--   then read out as 3456 fine channels.
----------------------------------------------------------------------------------
library IEEE, common_lib, filterbanks_lib;
use common_lib.common_pkg.all;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity correlatorFBTop25 is
    generic(
        METABITS : integer := 64;     -- Width in bits of the meta_i and meta_o ports.
        FRAMESTODROP : integer := 11  -- Number of output frames to drop after a reset (to account for initialisation of the filterbank)
    );
    port(
        -- clock, target is 380 MHz
        clk : in std_logic;
        rst : in std_logic;
        -- Data input, common valid signal, expects packets of 4096 samples. Requires at least 2 clocks idle time between packets.
        data0_i : in t_slv_8_arr(1 downto 0);  -- 4 Inputs, each complex data, 8 bit real, 8 bit imaginary.
        data1_i : in t_slv_8_arr(1 downto 0);
        data2_i : in t_slv_8_arr(1 downto 0);
        data3_i : in t_slv_8_arr(1 downto 0);
        meta_i  : in std_logic_vector((METABITS-1) downto 0);
        valid_i : in std_logic;
        -- Data out; bursts of 3456 clocks for each channel.
        data0_o : out t_slv_16_arr(1 downto 0);   -- 4 outputs, real and imaginary parts in (0) and (1) respectively;
        data1_o : out t_slv_16_arr(1 downto 0);
        data2_o : out t_slv_16_arr(1 downto 0);
        data3_o : out t_slv_16_arr(1 downto 0);
        meta_o  : out std_logic_vector((METABITS-1) downto 0);
        valid_o : out std_logic;
        -- Writing FIR Taps
        FIRTapData_i : in std_logic_vector(17 downto 0);  -- For register writes of the filtertaps.
        FIRTapData_o : out std_logic_vector(17 downto 0); -- For register reads of the filtertaps. 3 cycle latency from FIRTapAddr_i
        FIRTapAddr_i : in std_logic_vector(15 downto 0);  -- 4096 * 12 filter taps = 49152 total.
        FIRTapWE_i   : in std_logic;
        FIRTapClk    : in std_logic
    );
end correlatorFBTop25;

architecture Behavioral of correlatorFBTop25 is
    
    signal wrData64 : std_logic_vector(63 downto 0);
    signal FBmemRdData : t_slv_64_arr(11 downto 0);
    signal FBmemFIRTaps : t_slv_18_arr(11 downto 0);
    
    type fbtype is array(7 downto 0) of t_slv_8_arr(11 downto 0);
    signal FBRdData : fbtype; 
    signal FIRDout : t_slv_25_arr(7 downto 0);
    signal fftIndex : t_slv_12_arr(3 downto 0);
    
    signal fftRealOut : t_slv_16_arr(3 downto 0);
    signal fftImagOut : t_slv_16_arr(3 downto 0);
    signal fftvalidOut : std_logic_vector(3 downto 0) := "0000";
    
    signal startAdv : std_logic_vector(31 downto 0);
    signal validDel1, validDel2 : std_logic := '0';
    signal startFFT : std_logic := '0';
    
    signal reorderDout0, reorderDout1, reorderDout2, reorderDout3 : std_logic_vector(63 downto 0);
    signal reorderWE : std_logic_vector(1 downto 0);
    signal reorderWrAddr : std_logic_vector(11 downto 0);
    signal reorderRdAddr : std_logic_vector(11 downto 0);
    signal bufSelectWr, bufSelectRd : std_logic := '0';
    signal reorderDin0, reorderDin1 : std_logic_vector(63 downto 0);
    signal rdRunning : std_logic := '0';
    signal rdRunningDel2, rdRunningDel1 : std_logic := '0';
    signal validOutDel1 : std_logic := '0';
    signal bufSelectRdDel1, bufSelectRdDel2 : std_logic := '0';
    
    signal metaDel0, metaDel1, metaDel2, metaDel3, metaDel4 : std_logic_vector(METABITS+16-1 downto 0);
    signal metaOut : std_logic_vector((METABITS-1) downto 0);
    signal outputCountOut : std_logic_vector(15 downto 0);
    signal outputCount : std_logic_vector(15 downto 0);
    signal metaDel1Count, metaDel2Count, metaDel3Count : std_logic_vector(11 downto 0);
    
begin
    
    ------------------------------------------------------------------------------------
    -- 1. Input Memory
    -- ---------------
    
    wrData64 <= data3_i(1) & data3_i(0) & data2_i(1) & data2_i(0) & data1_i(1) & data1_i(0) & data0_i(1) & data0_i(0);

    cmem : entity filterbanks_lib.correlatorFBMem
    generic map (
        TAPS => 12)  -- Note only partially parameterized; modification needed to support anything other than 12.
    port map (
        clk      => clk,
        -- Write data for the start of the chain
        wrData_i => wrData64,         -- in(63:0);
        wrEn_i   => valid_i,          -- in std_logic; should be a burst of 4096 clocks.
        -- Read data, comes out 2 clocks after the first write.
        rd_data_o  => FBmemRdData,    -- out array64bit_type(TAPS-1 downto 0); -- 64 bits wide, 12 taps simultaneously; First sample is wr_data_i delayed by 1 clock. 
        coef_o     => FBmemFIRTaps,   -- out array18bit_type(TAPS-1 downto 0); -- 18 bits per filter tap.
        -- Writing FIR Taps
        FIRTapData_i => FIRTapData_i, -- in(17:0);  -- For register writes of the filtertaps.
        FIRTapData_o => FIRTapData_o, -- out(17:0); -- For register reads of the filtertaps. 3 cycle latency from FIRTapAddr_i
        FIRTapAddr_i => FIRTapAddr_i, -- in(15:0);  -- 4096 * 12 filter taps = 49152 total.
        FIRTapWE_i   => FIRTapWE_i,   -- in std_logic;
        FIRTapClk    => FIRTapClk     -- in std_logic
    );


    -------------------------------------------------------------------------------------
    -- 2. FIR filter
    -- -------------
    -- 8 instances, 4 channels * (real + imaginary). Same filter taps used for all.
    -- In low.CBF, processes simultaneously 2 (real+imaginary) * 2 (stations) * 2 (polarisations) = 8
    -- 
    
    CsampleGen : for j in 0 to 7 generate
        coefGen : for k in 0 to 11 generate
            FBRdData(j)(k) <= FBmemRdData(k)((j*8 + 7) downto (j*8));
        end generate;
    end generate;
    
    sampleGen : for j in 0 to 7 generate
            
        FIR : entity filterbanks_lib.fb_DSP25
        generic map (
            TAPS => 12)  -- The module instantiates this number of DSPs
        port map (
            clk    => clk,
            data_i => FBRdData(j),  -- in array8bit_type(11 downto 0);
            coef_i => FBmemFIRTaps, -- in array18bit_type(11 downto 0);
            data_o => FIRDout(j)    -- out(24:0)
        );
    
    end generate;
    
    -------------------------------------------------------------------------------------
    -- 3. FFT
    -- -----------------
    -- 4 x 4096 point FFTs.
    
    process(clk)
    begin
        if rising_edge(clk) then
            validDel1 <= valid_i;
            validDel2 <= validDel1;
            if validDel1 = '1' and validDel2 = '0' then
                startAdv(0) <= '1';
            else
                startAdv(0) <= '0';
            end if;
            
            startAdv(31 downto 1) <= startAdv(30 downto 0);
            startFFT <= startAdv(12); -- Delay accounts for the delay through the FIR filter 
            
            -- meta and output count
            -- Once a packet comes it data comes out after a fixed latency, but the gap between packets is variable.
            -- So we use a delay line which shifts after 4095 clocks if there is data in it. 
            if rst = '1' then
                outputCount <= (others => '0');
            elsif valid_i = '1' and validDel1 = '0' then -- rising edge of valid
                outputCount <= std_logic_vector(unsigned(outputCount) + 1);
                metaDel0 <= outputCount & meta_i;
            end if;
            
            if valid_i = '0' and validDel1 = '1' then -- falling edge of valid
                metaDel1 <= metaDel0;
                metaDel1Count <= "111111111111";
            elsif metaDel1Count /= "000000000000" then
                metaDel1Count <= std_logic_vector(unsigned(metaDel1Count) - 1);
            end if;
            
            if metaDel1Count = "000000000001" then
                metaDel2 <= metaDel1;
                metaDel2Count <= "111111111111";
            elsif metaDel2Count /= "000000000000" then
                metaDel2Count <= std_logic_vector(unsigned(metaDel2Count) - 1);
            end if;
            
            if metaDel2Count = "000000000001" then
                metaDel3 <= metaDel2;
                metaDel3Count <= "111111111111";
            elsif metaDel3Count /= "000000000000" then
                metaDel3Count <= std_logic_vector(unsigned(metaDel3Count) - 1);
            end if;
            
            if metaDel3Count = "000000000001" then
                metaDel4 <= metaDel3;
            end if;
            
            
        end if;
    end process;
    
    
    fftgen : for j in 0 to 3 generate
        
        fft4096 : entity filterbanks_lib.correlatorFFT25wrapper
        port map (
            clk  => clk,
            -- Input
            real_i  => FIRDout(j*2),     -- in(24:0); -- 25 bit real data
            imag_i  => FIRDout(j*2 + 1), -- in(24:0); -- 25 bit imaginary data
            start_i => startFFT,         -- in std_logic;                     -- pulse high; one clock in advance of the data ?
            -- Output
            real_o  => fftRealOut(j), -- out(15:0);
            imag_o  => fftImagOut(j), -- out(15:0);
            index_o => fftIndex(j),   -- out(11:0);
            valid_o => fftvalidOut(j) -- out std_logic
        );
    
    end generate;
    
    -------------------------------------------------------------------------------------
    -- 4. Reorder the output from bit-reversed to the central 3456 channels, low to high frequency. 
    -- 
    -- Uses an ultraRAM double buffer.
      
    process(clk)
    begin
        if rising_edge(clk) then
        
            if (fftvalidOut(0) = '1' and (signed(fftIndex(0)) > -1729) and (signed(fftIndex(0)) < 1728)) then
                if bufSelectWr = '0' then
                    reorderWE(0) <= '1';
                    reorderWE(1) <= '0';
                else
                    reorderWE(0) <= '0';
                    reorderWE(1) <= '1';
                end if;
            else
                reorderWE(0) <= '0';
                reorderWE(1) <= '0';
            end if;
            reorderWrAddr <= std_logic_vector(signed(fftIndex(0)) + 1728);
            reorderDin0 <= fftImagOut(1) & fftRealOut(1) & fftImagOut(0) & fftRealOut(0);
            reorderDin1 <= fftImagOut(3) & fftRealOut(3) & fftImagOut(2) & fftRealOut(2);
            
            -- Falling edge of validOut triggers reading of the data from the memory
            validOutDel1 <= fftvalidOut(0);
            if fftvalidOut(0) = '0' and validOutDel1 = '1' then
                reorderRdAddr <= "000000000000";
                bufSelectWr <= not bufSelectWr;
                bufSelectRd <= bufSelectWr;
                rdRunning <= '1';
            elsif rdRunning = '1' then
                reorderRdAddr <= std_logic_vector(unsigned(reorderRdAddr) + 1);
                -- read address runs from 0 to 3455
                if unsigned(reorderRdAddr) = 3455 then
                   rdRunning <= '0';
                end if;
            end if;
            rdRunningDel1 <= rdRunning;
            rdRunningDel2 <= rdRunningDel1;
            bufSelectRdDel1 <= bufSelectRd;
            bufSelectRdDel2 <= bufSelectRdDel1;
        end if;
    end process;

    -- Two URAMs for first half of the double buffer
    reorderURAM0 : entity filterbanks_lib.URAMWrapper
    port map (
        clk => clk,
        -- write side
        wrAddr => reorderWrAddr, -- in(11:0);
        din    => reorderDin0,   -- in(63:0);
        we     => reorderWE(0),  -- in std_logic;
        -- read side
        rdAddr => reorderRdAddr, -- in(11:0);
        dout   => reorderDout0   -- out(63:0)
    );

    reorderURAM1 : entity filterbanks_lib.URAMWrapper
    port map (
        clk => clk,
        -- write side
        wrAddr => reorderWrAddr, -- in(11:0);
        din    => reorderDin1,   -- in(63:0);
        we     => reorderWE(0),  -- in std_logic;
        -- read side
        rdAddr => reorderRdAddr, -- in(11:0);
        dout   => reorderDout1   -- out(63:0)
    );    
    
    -- Two URAMs for the second half of the double buffer
    reorderURAM2 : entity filterbanks_lib.URAMWrapper
    port map (
        clk => clk,
        -- write side
        wrAddr => reorderWrAddr, -- in(11:0);
        din    => reorderDin0,   -- in(63:0);
        we     => reorderWE(1),  -- in std_logic;
        -- read side
        rdAddr => reorderRdAddr, -- in(11:0);
        dout   => reorderDout2   -- out(63:0)
    );

    reorderURAM3 : entity filterbanks_lib.URAMWrapper
    port map (
        clk => clk,
        -- write side
        wrAddr => reorderWrAddr, -- in(11:0);
        din    => reorderDin1,   -- in(63:0);
        we     => reorderWE(1),  -- in std_logic;
        -- read side
        rdAddr => reorderRdAddr, -- in(11:0);
        dout   => reorderDout3   -- out(63:0)
    );    
    

    process(clk)
    begin
        if rising_edge(clk) then
            if rdRunningDel1 = '1' and rdRunningDel2 = '0' then -- Rising edge of rdRunning, two clocks prior to valid_o
                metaOut <= metaDel2((METABITS-1) downto 0);
                outputCountOut <= metaDel2((METABITS+15) downto METABITS);
            end if;
            
            if bufSelectRdDel2 = '0' then
                data0_o(0) <= reorderDout0(15 downto 0);
                data0_o(1) <= reorderDout0(31 downto 16);
                data1_o(0) <= reorderDout0(47 downto 32);
                data1_o(1) <= reorderDout0(63 downto 48);
                data2_o(0) <= reorderDout1(15 downto 0);
                data2_o(1) <= reorderDout1(31 downto 16);
                data3_o(0) <= reorderDout1(47 downto 32);
                data3_o(1) <= reorderDout1(63 downto 48);
            else
                data0_o(0) <= reorderDout2(15 downto 0);
                data0_o(1) <= reorderDout2(31 downto 16);
                data1_o(0) <= reorderDout2(47 downto 32);
                data1_o(1) <= reorderDout2(63 downto 48);
                data2_o(0) <= reorderDout3(15 downto 0);
                data2_o(1) <= reorderDout3(31 downto 16);
                data3_o(0) <= reorderDout3(47 downto 32);
                data3_o(1) <= reorderDout3(63 downto 48);
            end if;
            
            if (unsigned(outputCountOut) >= FRAMESTODROP) then
                valid_o <= rdRunningDel2;
            else
                valid_o <= '0';
            end if;
            
        end if;
    end process;    
    
    meta_o <= metaOut;
    
end Behavioral;
