
// file: ibert_bank_gth.v
//////////////////////////////////////////////////////////////////////////////
//   ____  ____ 
//  /   /\/   /
// /___/  \  /    Vendor: Xilinx
// \   \   \/     Version : 2012.3
//  \   \         Application : IBERT 7Series 
//  /   /         Filename : example_ibert_bank_gth
// /___/   /\     
// \   \  /  \ 
//  \___\/\___\
//
//
// Module example_ibert_bank_gth
// Generated by Xilinx IBERT_7S 
//////////////////////////////////////////////////////////////////////////////

`define C_NUM_GTH_QUADS 13
`define C_GTH_REFCLKS_USED 6
module example_ibert_bank_gth
(
  // GT top level ports
  output [(4*`C_NUM_GTH_QUADS)-1:0]		gth_txn_o,
  output [(4*`C_NUM_GTH_QUADS)-1:0]		gth_txp_o,
  input  [(4*`C_NUM_GTH_QUADS)-1:0]    	gth_rxn_i,
  input  [(4*`C_NUM_GTH_QUADS)-1:0]   	gth_rxp_i,
  input                           	gth_sysclkp_i,
  input                           	gth_sysclkn_i,
  input  [`C_GTH_REFCLKS_USED-1:0]      gth_refclk0p_i,
  input  [`C_GTH_REFCLKS_USED-1:0]      gth_refclk0n_i,
  input  [`C_GTH_REFCLKS_USED-1:0]      gth_refclk1p_i,
  input  [`C_GTH_REFCLKS_USED-1:0]      gth_refclk1n_i,
  input [0:0]ferr_n_tri_i,
  output [0:0]hmc_refclk_sel_tri_o,
  inout iic_main_scl_io,
  inout iic_main_sda_io,
  output [2:0]iic_mux_reset_b,
  output [1:0]lxrxps_tri_o,
  input [1:0]lxtxps_tri_i,
  output [1:0]refclk_boot_tri_o,
  input reset,
  input rs232_uart_rxd,
  output rs232_uart_txd
);

  //
  // Ibert refclk internal signals
  //
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk0_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk1_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk0_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk1_i;        	
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk0_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk1_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk00_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk10_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk01_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qrefclk11_i;  
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk00_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk10_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk01_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qnorthrefclk11_i;  
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk00_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk10_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk01_i;
  wire  [`C_NUM_GTH_QUADS-1:0]    gth_qsouthrefclk11_i; 
  wire  [`C_GTH_REFCLKS_USED-1:0] gth_refclk0_i;
  wire  [`C_GTH_REFCLKS_USED-1:0] gth_refclk1_i;
  wire  [`C_GTH_REFCLKS_USED-1:0] gth_odiv2_0_i;
  wire  [`C_GTH_REFCLKS_USED-1:0] gth_odiv2_1_i;
  wire                        gth_sysclk_i;
  wire [0:0]ferr_n_tri_i;
  wire [0:0]hmc_refclk_sel_tri_o;
  wire iic_main_scl_i;
  wire iic_main_scl_io;
  wire iic_main_scl_o;
  wire iic_main_scl_t;
  wire iic_main_sda_i;
  wire iic_main_sda_io;
  wire iic_main_sda_o;
  wire iic_main_sda_t;
  wire [2:0]iic_mux_reset_b;
  wire [1:0]lxrxps_tri_o;
  wire [1:0]lxtxps_tri_i;
  wire [1:0]refclk_boot_tri_o;
  wire reset;
  wire rs232_uart_rxd;
  wire rs232_uart_txd;

  //
  // Refclk IBUFDS instantiations
  //
    IBUFDS_GTE3 u_buf_gth_q2_clk0
      (
        .O            (gth_refclk0_i[0]),
        .ODIV2        (gth_odiv2_0_i[0]),
        .CEB          (1'b0),
        .I            (gth_refclk0p_i[0]),
        .IB           (gth_refclk0n_i[0])
      );

    IBUFDS_GTE3 u_buf_gth_q2_clk1
      (
        .O            (gth_refclk1_i[0]),
        .ODIV2        (gth_odiv2_1_i[0]),
        .CEB          (1'b0),
        .I            (gth_refclk1p_i[0]),
        .IB           (gth_refclk1n_i[0])
      );
    IBUFDS_GTE3 u_buf_gth_q3_clk0
      (
        .O            (gth_refclk0_i[1]),
        .ODIV2        (gth_odiv2_0_i[1]),
        .CEB          (1'b0),
        .I            (gth_refclk0p_i[1]),
        .IB           (gth_refclk0n_i[1])
      );

    IBUFDS_GTE3 u_buf_gth_q3_clk1
      (
        .O            (gth_refclk1_i[1]),
        .ODIV2        (gth_odiv2_1_i[1]),
        .CEB          (1'b0),
        .I            (gth_refclk1p_i[1]),
        .IB           (gth_refclk1n_i[1])
      );
    IBUFDS_GTE3 u_buf_gth_q5_clk0
      (
        .O            (gth_refclk0_i[2]),
        .ODIV2        (gth_odiv2_0_i[2]),
        .CEB          (1'b0),
        .I            (gth_refclk0p_i[2]),
        .IB           (gth_refclk0n_i[2])
      );

    IBUFDS_GTE3 u_buf_gth_q5_clk1
      (
        .O            (gth_refclk1_i[2]),
        .ODIV2        (gth_odiv2_1_i[2]),
        .CEB          (1'b0),
        .I            (gth_refclk1p_i[2]),
        .IB           (gth_refclk1n_i[2])
      );
    IBUFDS_GTE3 u_buf_gth_q7_clk0
      (
        .O            (gth_refclk0_i[3]),
        .ODIV2        (gth_odiv2_0_i[3]),
        .CEB          (1'b0),
        .I            (gth_refclk0p_i[3]),
        .IB           (gth_refclk0n_i[3])
      );

    IBUFDS_GTE3 u_buf_gth_q7_clk1
      (
        .O            (gth_refclk1_i[3]),
        .ODIV2        (gth_odiv2_1_i[3]),
        .CEB          (1'b0),
        .I            (gth_refclk1p_i[3]),
        .IB           (gth_refclk1n_i[3])
      );
    IBUFDS_GTE3 u_buf_gth_q11_clk0
      (
        .O            (gth_refclk0_i[4]),
        .ODIV2        (gth_odiv2_0_i[4]),
        .CEB          (1'b0),
        .I            (gth_refclk0p_i[4]),
        .IB           (gth_refclk0n_i[4])
      );

    IBUFDS_GTE3 u_buf_gth_q11_clk1
      (
        .O            (gth_refclk1_i[4]),
        .ODIV2        (gth_odiv2_1_i[4]),
        .CEB          (1'b0),
        .I            (gth_refclk1p_i[4]),
        .IB           (gth_refclk1n_i[4])
      );
    IBUFDS_GTE3 u_buf_gth_q14_clk0
      (
        .O            (gth_refclk0_i[5]),
        .ODIV2        (gth_odiv2_0_i[5]),
        .CEB          (1'b0),
        .I            (gth_refclk0p_i[5]),
        .IB           (gth_refclk0n_i[5])
      );

    IBUFDS_GTE3 u_buf_gth_q14_clk1
      (
        .O            (gth_refclk1_i[5]),
        .ODIV2        (gth_odiv2_1_i[5]),
        .CEB          (1'b0),
        .I            (gth_refclk1p_i[5]),
        .IB           (gth_refclk1n_i[5])
      );

  //
  // Refclk connection from each IBUFDS to respective quads depending on the source selected in gui
  //
  assign gth_qrefclk0_i[0] = 1'b0;
  assign gth_qrefclk1_i[0] = 1'b0;
  assign gth_qnorthrefclk0_i[0] = 1'b0;
  assign gth_qnorthrefclk1_i[0] = 1'b0;
  assign gth_qsouthrefclk0_i[0] = gth_refclk0_i[0];
  assign gth_qsouthrefclk1_i[0] = 1'b0;
//COMMON clock connection
  assign gth_qrefclk00_i[0] = 1'b0;
  assign gth_qrefclk10_i[0] = 1'b0;
  assign gth_qrefclk01_i[0] = 1'b0;
  assign gth_qrefclk11_i[0] = 1'b0;
  assign gth_qnorthrefclk00_i[0] = 1'b0;
  assign gth_qnorthrefclk10_i[0] = 1'b0;
  assign gth_qnorthrefclk01_i[0] = 1'b0;
  assign gth_qnorthrefclk11_i[0] = 1'b0;
  assign gth_qsouthrefclk00_i[0] = gth_refclk0_i[0];
  assign gth_qsouthrefclk10_i[0] = 1'b0;
  assign gth_qsouthrefclk01_i[0] = 1'b0;
  assign gth_qsouthrefclk11_i[0] = 1'b0;
 
  assign gth_qrefclk0_i[1] = gth_refclk0_i[0];
  assign gth_qrefclk1_i[1] = gth_refclk1_i[0];
  assign gth_qnorthrefclk0_i[1] = 1'b0;
  assign gth_qnorthrefclk1_i[1] = 1'b0;
  assign gth_qsouthrefclk0_i[1] = 1'b0;
  assign gth_qsouthrefclk1_i[1] = 1'b0;
//COMMON clock connection
  assign gth_qrefclk00_i[1] = gth_refclk0_i[0];
  assign gth_qrefclk10_i[1] = gth_refclk1_i[0];
  assign gth_qrefclk01_i[1] = 1'b0;
  assign gth_qrefclk11_i[1] = 1'b0;  
  assign gth_qnorthrefclk00_i[1] = 1'b0;
  assign gth_qnorthrefclk10_i[1] = 1'b0;
  assign gth_qnorthrefclk01_i[1] = 1'b0;
  assign gth_qnorthrefclk11_i[1] = 1'b0;  
  assign gth_qsouthrefclk00_i[1] = 1'b0;
  assign gth_qsouthrefclk10_i[1] = 1'b0;  
  assign gth_qsouthrefclk01_i[1] = 1'b0;
  assign gth_qsouthrefclk11_i[1] = 1'b0; 
 

  assign gth_qrefclk0_i[2] = gth_refclk0_i[1];
  assign gth_qrefclk1_i[2] = gth_refclk1_i[1];
  assign gth_qnorthrefclk0_i[2] = 1'b0;
  assign gth_qnorthrefclk1_i[2] = 1'b0;
  assign gth_qsouthrefclk0_i[2] = 1'b0;
  assign gth_qsouthrefclk1_i[2] = 1'b0;
//COMMON clock connection
  assign gth_qrefclk00_i[2] = gth_refclk0_i[1];
  assign gth_qrefclk10_i[2] = gth_refclk1_i[1];
  assign gth_qrefclk01_i[2] = 1'b0;
  assign gth_qrefclk11_i[2] = 1'b0;  
  assign gth_qnorthrefclk00_i[2] = 1'b0;
  assign gth_qnorthrefclk10_i[2] = 1'b0;
  assign gth_qnorthrefclk01_i[2] = 1'b0;
  assign gth_qnorthrefclk11_i[2] = 1'b0;  
  assign gth_qsouthrefclk00_i[2] = 1'b0;
  assign gth_qsouthrefclk10_i[2] = 1'b0;  
  assign gth_qsouthrefclk01_i[2] = 1'b0;
  assign gth_qsouthrefclk11_i[2] = 1'b0; 
 

  assign gth_qrefclk0_i[3] = gth_refclk0_i[2];
  assign gth_qrefclk1_i[3] = gth_refclk1_i[2];
  assign gth_qnorthrefclk0_i[3] = 1'b0;
  assign gth_qnorthrefclk1_i[3] = 1'b0;
  assign gth_qsouthrefclk0_i[3] = 1'b0;
  assign gth_qsouthrefclk1_i[3] = 1'b0;
//COMMON clock connection
  assign gth_qrefclk00_i[3] = gth_refclk0_i[2];
  assign gth_qrefclk10_i[3] = gth_refclk1_i[2];
  assign gth_qrefclk01_i[3] = 1'b0;
  assign gth_qrefclk11_i[3] = 1'b0;  
  assign gth_qnorthrefclk00_i[3] = 1'b0;
  assign gth_qnorthrefclk10_i[3] = 1'b0;
  assign gth_qnorthrefclk01_i[3] = 1'b0;
  assign gth_qnorthrefclk11_i[3] = 1'b0;  
  assign gth_qsouthrefclk00_i[3] = 1'b0;
  assign gth_qsouthrefclk10_i[3] = 1'b0;  
  assign gth_qsouthrefclk01_i[3] = 1'b0;
  assign gth_qsouthrefclk11_i[3] = 1'b0; 
 

  assign gth_qrefclk0_i[4] = 1'b0;
  assign gth_qrefclk1_i[4] = 1'b0;
  assign gth_qnorthrefclk0_i[4] = 1'b0;
  assign gth_qnorthrefclk1_i[4] = 1'b0;
  assign gth_qsouthrefclk0_i[4] = gth_refclk0_i[3];
  assign gth_qsouthrefclk1_i[4] = 1'b0;
//COMMON clock connection
  assign gth_qrefclk00_i[4] = 1'b0;
  assign gth_qrefclk10_i[4] = 1'b0;
  assign gth_qrefclk01_i[4] = 1'b0;
  assign gth_qrefclk11_i[4] = 1'b0;
  assign gth_qnorthrefclk00_i[4] = 1'b0;
  assign gth_qnorthrefclk10_i[4] = 1'b0;
  assign gth_qnorthrefclk01_i[4] = 1'b0;
  assign gth_qnorthrefclk11_i[4] = 1'b0;
  assign gth_qsouthrefclk00_i[4] = gth_refclk0_i[3];
  assign gth_qsouthrefclk10_i[4] = 1'b0;
  assign gth_qsouthrefclk01_i[4] = 1'b0;
  assign gth_qsouthrefclk11_i[4] = 1'b0;
 
  assign gth_qrefclk0_i[5] = gth_refclk0_i[3];
  assign gth_qrefclk1_i[5] = gth_refclk1_i[3];
  assign gth_qnorthrefclk0_i[5] = 1'b0;
  assign gth_qnorthrefclk1_i[5] = 1'b0;
  assign gth_qsouthrefclk0_i[5] = 1'b0;
  assign gth_qsouthrefclk1_i[5] = 1'b0;
//COMMON clock connection
  assign gth_qrefclk00_i[5] = gth_refclk0_i[3];
  assign gth_qrefclk10_i[5] = gth_refclk1_i[3];
  assign gth_qrefclk01_i[5] = 1'b0;
  assign gth_qrefclk11_i[5] = 1'b0;  
  assign gth_qnorthrefclk00_i[5] = 1'b0;
  assign gth_qnorthrefclk10_i[5] = 1'b0;
  assign gth_qnorthrefclk01_i[5] = 1'b0;
  assign gth_qnorthrefclk11_i[5] = 1'b0;  
  assign gth_qsouthrefclk00_i[5] = 1'b0;
  assign gth_qsouthrefclk10_i[5] = 1'b0;  
  assign gth_qsouthrefclk01_i[5] = 1'b0;
  assign gth_qsouthrefclk11_i[5] = 1'b0; 
 

  assign gth_qrefclk0_i[6] = 1'b0;
  assign gth_qrefclk1_i[6] = 1'b0;
  assign gth_qnorthrefclk0_i[6] = gth_refclk0_i[3];
  assign gth_qnorthrefclk1_i[6] = 1'b0;
  assign gth_qsouthrefclk0_i[6] = 1'b0;
  assign gth_qsouthrefclk1_i[6] = 1'b0;
//COMMON clock connection
  assign gth_qrefclk00_i[6] = 1'b0;
  assign gth_qrefclk10_i[6] = 1'b0;
  assign gth_qrefclk01_i[6] = 1'b0;
  assign gth_qrefclk11_i[6] = 1'b0;
  assign gth_qnorthrefclk00_i[6] = gth_refclk0_i[3];
  assign gth_qnorthrefclk10_i[6] = 1'b0;
  assign gth_qnorthrefclk01_i[6] = 1'b0;
  assign gth_qnorthrefclk11_i[6] = 1'b0;
  assign gth_qsouthrefclk00_i[6] = 1'b0;
  assign gth_qsouthrefclk10_i[6] = 1'b0;
  assign gth_qsouthrefclk01_i[6] = 1'b0;
  assign gth_qsouthrefclk11_i[6] = 1'b0;
 
  assign gth_qrefclk0_i[7] = 1'b0;
  assign gth_qrefclk1_i[7] = 1'b0;
  assign gth_qnorthrefclk0_i[7] = gth_refclk0_i[3];
  assign gth_qnorthrefclk1_i[7] = 1'b0;
  assign gth_qsouthrefclk0_i[7] = 1'b0;
  assign gth_qsouthrefclk1_i[7] = 1'b0;
//COMMON clock connection
  assign gth_qrefclk00_i[7] = 1'b0;
  assign gth_qrefclk10_i[7] = 1'b0;
  assign gth_qrefclk01_i[7] = 1'b0;
  assign gth_qrefclk11_i[7] = 1'b0;
  assign gth_qnorthrefclk00_i[7] = gth_refclk0_i[3];
  assign gth_qnorthrefclk10_i[7] = 1'b0;
  assign gth_qnorthrefclk01_i[7] = 1'b0;
  assign gth_qnorthrefclk11_i[7] = 1'b0;
  assign gth_qsouthrefclk00_i[7] = 1'b0;
  assign gth_qsouthrefclk10_i[7] = 1'b0;
  assign gth_qsouthrefclk01_i[7] = 1'b0;
  assign gth_qsouthrefclk11_i[7] = 1'b0;
 
  assign gth_qrefclk0_i[8] = 1'b0;
  assign gth_qrefclk1_i[8] = 1'b0;
  assign gth_qnorthrefclk0_i[8] = 1'b0;
  assign gth_qnorthrefclk1_i[8] = 1'b0;
  assign gth_qsouthrefclk0_i[8] = gth_refclk0_i[4];
  assign gth_qsouthrefclk1_i[8] = 1'b0;
//COMMON clock connection
  assign gth_qrefclk00_i[8] = 1'b0;
  assign gth_qrefclk10_i[8] = 1'b0;
  assign gth_qrefclk01_i[8] = 1'b0;
  assign gth_qrefclk11_i[8] = 1'b0;
  assign gth_qnorthrefclk00_i[8] = 1'b0;
  assign gth_qnorthrefclk10_i[8] = 1'b0;
  assign gth_qnorthrefclk01_i[8] = 1'b0;
  assign gth_qnorthrefclk11_i[8] = 1'b0;
  assign gth_qsouthrefclk00_i[8] = gth_refclk0_i[4];
  assign gth_qsouthrefclk10_i[8] = 1'b0;
  assign gth_qsouthrefclk01_i[8] = 1'b0;
  assign gth_qsouthrefclk11_i[8] = 1'b0;
 
  assign gth_qrefclk0_i[9] = gth_refclk0_i[4];
  assign gth_qrefclk1_i[9] = gth_refclk1_i[4];
  assign gth_qnorthrefclk0_i[9] = 1'b0;
  assign gth_qnorthrefclk1_i[9] = 1'b0;
  assign gth_qsouthrefclk0_i[9] = 1'b0;
  assign gth_qsouthrefclk1_i[9] = 1'b0;
//COMMON clock connection
  assign gth_qrefclk00_i[9] = gth_refclk0_i[4];
  assign gth_qrefclk10_i[9] = gth_refclk1_i[4];
  assign gth_qrefclk01_i[9] = 1'b0;
  assign gth_qrefclk11_i[9] = 1'b0;  
  assign gth_qnorthrefclk00_i[9] = 1'b0;
  assign gth_qnorthrefclk10_i[9] = 1'b0;
  assign gth_qnorthrefclk01_i[9] = 1'b0;
  assign gth_qnorthrefclk11_i[9] = 1'b0;  
  assign gth_qsouthrefclk00_i[9] = 1'b0;
  assign gth_qsouthrefclk10_i[9] = 1'b0;  
  assign gth_qsouthrefclk01_i[9] = 1'b0;
  assign gth_qsouthrefclk11_i[9] = 1'b0; 
 

  assign gth_qrefclk0_i[10] = 1'b0;
  assign gth_qrefclk1_i[10] = 1'b0;
  assign gth_qnorthrefclk0_i[10] = gth_refclk0_i[4];
  assign gth_qnorthrefclk1_i[10] = 1'b0;
  assign gth_qsouthrefclk0_i[10] = 1'b0;
  assign gth_qsouthrefclk1_i[10] = 1'b0;
//COMMON clock connection
  assign gth_qrefclk00_i[10] = 1'b0;
  assign gth_qrefclk10_i[10] = 1'b0;
  assign gth_qrefclk01_i[10] = 1'b0;
  assign gth_qrefclk11_i[10] = 1'b0;
  assign gth_qnorthrefclk00_i[10] = gth_refclk0_i[4];
  assign gth_qnorthrefclk10_i[10] = 1'b0;
  assign gth_qnorthrefclk01_i[10] = 1'b0;
  assign gth_qnorthrefclk11_i[10] = 1'b0;
  assign gth_qsouthrefclk00_i[10] = 1'b0;
  assign gth_qsouthrefclk10_i[10] = 1'b0;
  assign gth_qsouthrefclk01_i[10] = 1'b0;
  assign gth_qsouthrefclk11_i[10] = 1'b0;
 
  assign gth_qrefclk0_i[11] = 1'b0;
  assign gth_qrefclk1_i[11] = 1'b0;
  assign gth_qnorthrefclk0_i[11] = gth_refclk0_i[4];
  assign gth_qnorthrefclk1_i[11] = 1'b0;
  assign gth_qsouthrefclk0_i[11] = 1'b0;
  assign gth_qsouthrefclk1_i[11] = 1'b0;
//COMMON clock connection
  assign gth_qrefclk00_i[11] = 1'b0;
  assign gth_qrefclk10_i[11] = 1'b0;
  assign gth_qrefclk01_i[11] = 1'b0;
  assign gth_qrefclk11_i[11] = 1'b0;
  assign gth_qnorthrefclk00_i[11] = gth_refclk0_i[4];
  assign gth_qnorthrefclk10_i[11] = 1'b0;
  assign gth_qnorthrefclk01_i[11] = 1'b0;
  assign gth_qnorthrefclk11_i[11] = 1'b0;
  assign gth_qsouthrefclk00_i[11] = 1'b0;
  assign gth_qsouthrefclk10_i[11] = 1'b0;
  assign gth_qsouthrefclk01_i[11] = 1'b0;
  assign gth_qsouthrefclk11_i[11] = 1'b0;
 
  assign gth_qrefclk0_i[12] = gth_refclk0_i[5];
  assign gth_qrefclk1_i[12] = gth_refclk1_i[5];
  assign gth_qnorthrefclk0_i[12] = 1'b0;
  assign gth_qnorthrefclk1_i[12] = 1'b0;
  assign gth_qsouthrefclk0_i[12] = 1'b0;
  assign gth_qsouthrefclk1_i[12] = 1'b0;
//COMMON clock connection
  assign gth_qrefclk00_i[12] = gth_refclk0_i[5];
  assign gth_qrefclk10_i[12] = gth_refclk1_i[5];
  assign gth_qrefclk01_i[12] = 1'b0;
  assign gth_qrefclk11_i[12] = 1'b0;  
  assign gth_qnorthrefclk00_i[12] = 1'b0;
  assign gth_qnorthrefclk10_i[12] = 1'b0;
  assign gth_qnorthrefclk01_i[12] = 1'b0;
  assign gth_qnorthrefclk11_i[12] = 1'b0;  
  assign gth_qsouthrefclk00_i[12] = 1'b0;
  assign gth_qsouthrefclk10_i[12] = 1'b0;  
  assign gth_qsouthrefclk01_i[12] = 1'b0;
  assign gth_qsouthrefclk11_i[12] = 1'b0; 
 

  //
  // Sysclock IBUFDS instantiation
  //
  IBUFGDS 
   #(.DIFF_TERM("FALSE"))
   u_ibufgds
    (
      .I(gth_sysclkp_i),
      .IB(gth_sysclkn_i),
      .O(gth_sysclk_i)
    );


  //
  // IBERT core instantiation
  //
  ibert_bank_gth u_ibert_gth_core
    (
      .txn_o(gth_txn_o),
      .txp_o(gth_txp_o),
      .rxn_i(gth_rxn_i),
      .rxp_i(gth_rxp_i),
      .clk(gth_sysclk_i),
      .gtrefclk0_i(gth_qrefclk0_i),
      .gtrefclk1_i(gth_qrefclk1_i),
      .gtnorthrefclk0_i(gth_qnorthrefclk0_i),
      .gtnorthrefclk1_i(gth_qnorthrefclk1_i),
      .gtsouthrefclk0_i(gth_qsouthrefclk0_i),
      .gtsouthrefclk1_i(gth_qsouthrefclk1_i),
      .gtrefclk00_i(gth_qrefclk00_i),
      .gtrefclk10_i(gth_qrefclk10_i),
      .gtrefclk01_i(gth_qrefclk01_i),
      .gtrefclk11_i(gth_qrefclk11_i),
      .gtnorthrefclk00_i(gth_qnorthrefclk00_i),
      .gtnorthrefclk10_i(gth_qnorthrefclk10_i),
      .gtnorthrefclk01_i(gth_qnorthrefclk01_i),
      .gtnorthrefclk11_i(gth_qnorthrefclk11_i),
      .gtsouthrefclk00_i(gth_qsouthrefclk00_i),
      .gtsouthrefclk10_i(gth_qsouthrefclk10_i),
      .gtsouthrefclk01_i(gth_qsouthrefclk01_i),
      .gtsouthrefclk11_i(gth_qsouthrefclk11_i)
    );

  IOBUF iic_main_scl_iobuf
       (.I(iic_main_scl_o),
        .IO(iic_main_scl_io),
        .O(iic_main_scl_i),
        .T(iic_main_scl_t));
  IOBUF iic_main_sda_iobuf
       (.I(iic_main_sda_o),
        .IO(iic_main_sda_io),
        .O(iic_main_sda_i),
        .T(iic_main_sda_t));
  system system_i
       (.FERR_N_tri_i(ferr_n_tri_i),
        .HMC_REFCLK_SEL_tri_o(hmc_refclk_sel_tri_o),
        .LxRXPS_tri_o(lxrxps_tri_o),
        .LxTXPS_tri_i(lxtxps_tri_i),
        .REFCLK_BOOT_tri_o(refclk_boot_tri_o),
        .gth_sysclk_i(gth_sysclk_i),
        .iic_main_scl_i(iic_main_scl_i),
        .iic_main_scl_o(iic_main_scl_o),
        .iic_main_scl_t(iic_main_scl_t),
        .iic_main_sda_i(iic_main_sda_i),
        .iic_main_sda_o(iic_main_sda_o),
        .iic_main_sda_t(iic_main_sda_t),
        .iic_mux_reset_b(iic_mux_reset_b),
        .reset(reset),
        .rs232_uart_rxd(rs232_uart_rxd),
        .rs232_uart_txd(rs232_uart_txd));

endmodule
