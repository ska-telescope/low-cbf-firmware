----------------------------------------------------------------------------------
-- Company: CSIRO CASS 
-- Engineer: David Humphrey
-- 
-- Create Date: 14.11.2018 11:27:29
-- Module Name: PSSFBTop - Behavioral
-- Description: 
--  Filterbank with 12 FIR taps, 64 point FFT, critically sampled.
--  Designed for the low.CBF PSS beamformer. Output is the central 54 frequency channels.
--  Processes 6 parallel signals, each with 8 bit complex data (8 bit real + 8 bit imaginary).
--  
-- Supporting Code:
--  The Matlab model should be in the directory ../matlab_model
--  Key files:
--   * ../matlab_model/run_PSSFB.m 
--       Generates input files for the simulation, runs the matlab model and compares with simulation output.
--   * ../matlab_model/get_rom_coefficients.m
--       Generates ROM data used in the firmware. ROMs are initialised using .coe files.
--       "PSSFIRTapsX.coe" : X runs from 1 to 12, contents of the 12 ROMS used to store the FIR filter taps.
--
--  Supporting VHDL 
--   * PSSFBtesttop.vhd 
--      Top level module that can be used to build this in a standalone version.
--   * PSSFB_tb.vhd
--      testbench, reads input data generated by the matlab code, and generates output data in text files for analysis by the matlab code. 
--
-- Structure:
--
--  File Structure
--  --------------
--  Outline of the structure shown below. Excludes most .xci files for DSPs, RAMs and ROMs.
--
--    PSSFBTop.vhd : This file, 6 complex inputs, 12 FIR filter taps, 64 point FFT, critically sampled
--        |
--        +-- PSSFBmem.vhd   : Input memory for the filterbank, 12 blocks of memory chained together, see "step 1. Filterbank memory" below.
--        +-- fb_DSP.vhd     : 12 TAP FIR filter, see "2. FIR filter" below.
--        +-- PSSFFTwrapper.vhd : 64 point FFT. see "3. 1280 point FFT" below.
--                |
--                +-- fft64_16bit.xci : standard Xilinx 64 point FFT
--
--  Resource Use
--  ------------
--  Approximate resource usage is 
--   LUTs = 7941
--   DSPs = 192
--   Registers = 13804
--   BRAMs (36K) = 9
--
--  Power (estimate based on related measurements on the zcu111 board)
--   about 1 W static, 3.5 W dynamic.
--   
--  -----------------------------------------------------------------------------------------------
--  Description
--  -----------
--
-- 1. Filterbank Memory
--   The filterbank memory consists of 11 blocks of memory chained together.
--   The read data from each memory is used both by the FIR filter and to write to the next memory in the chain.
--   The read and write addresses are staggered by one clock for each memory, implemented as a 12 sample delay line on
--   the address. This makes the timing easy to meet for the  memory address signals (which would otherwise be high-fanout signals)
--   and also enables use of the adders in the DSPs for the FIR filter.  
--
-- 2. FIR filter
--   The FIR filter uses 12 DSPs for each of the 12 simultaneous samples (6 channels * 2 (re+im)) that are read from the memory.
--   So the FIR filter uses (12 DSPS) * (6 simultaneous samples) * (2 (re+im)) = 144 DSPs.
--   The filter is implemented entirely in DSPs. The PCOUT port on the DSP is used to send the result of the multiplication
--   to the next DSP in the chain, where it is added using the adder in the DSP. This scheme requires that the inputs to the
--   12 DSPs are staggered to account for the pipeline stage on the PCOUT port. The staggering is done by controlling the address
--   to the memories as described above.
--
-- 3. 64 point FFT
--   Standard Xilinx FFT. Some messy logic at the front to account for the delay inserted by the "real-time" mode.
-- 
-- 4. Reorder memory
--   Data out of the FFT is in bit reversed order. It is stored in a double buffer in order from low to high frequencies,
--   then read out as 54 fine channels.
----------------------------------------------------------------------------------
library IEEE, common_lib, filterbanks_lib;
use IEEE.STD_LOGIC_1164.ALL;
use common_lib.common_pkg.all;
use IEEE.NUMERIC_STD.ALL;

entity PSSFBTop is
    port(
        -- clock, target is 380 MHz
        clk         : in std_logic;
        rst         : in std_logic;
        FIRTapUse_i : in std_logic;   -- FIR Taps are double buffered, choose which set of TAPs to use.
        -- Data input, common valid signal, expects packets of 64 samples. Requires at least 2 clocks idle time between packets.
        data0_i : in t_slv_8_arr(1 downto 0);  -- 6 Inputs, each complex data, 8 bit real, 8 bit imaginary.
        data1_i : in t_slv_8_arr(1 downto 0);
        data2_i : in t_slv_8_arr(1 downto 0);
        data3_i : in t_slv_8_arr(1 downto 0);
        data4_i : in t_slv_8_arr(1 downto 0);
        data5_i : in t_slv_8_arr(1 downto 0);
        valid_i : in std_logic;
        -- Data out; bursts of 54 clocks for each channel.
        data0_o : out t_slv_16_arr(1 downto 0);   -- 6 outputs, real and imaginary parts in (0) and (1) respectively;
        data1_o : out t_slv_16_arr(1 downto 0);
        data2_o : out t_slv_16_arr(1 downto 0);
        data3_o : out t_slv_16_arr(1 downto 0);
        data4_o : out t_slv_16_arr(1 downto 0);
        data5_o : out t_slv_16_arr(1 downto 0);
        valid_o : out std_logic;
        -- Writing FIR Taps
        FIRTapData_i   : in std_logic_vector(17 downto 0);  -- For register writes of the filtertaps.
        FIRTapData_o   : out std_logic_vector(17 downto 0); -- For register reads of the filtertaps. 3 cycle latency from FIRTapAddr_i
        FIRTapAddr_i   : in std_logic_vector(9 downto 0);   -- 64 * 12 filter taps = 768 total.
        FIRTapWE_i     : in std_logic;
        FIRTapClk      : in std_logic;
        FIRTapSelect_i : in std_logic  -- FIR Taps are double buffered; This selects the buffer to access for registers. Choose which buffer to use with FIRTapUse_i
    );
end PSSFBTop;

architecture Behavioral of PSSFBTop is

    -- reorder memory
    -- 1.5 BRAMs, simple dual port, 2 cycle read latency.
    -- Tcl:
    --  create_ip -name blk_mem_gen -vendor xilinx.com -library ip -version 8.4 -module_name PSSFBReorderMem -dir C:/projects/perentie/xilinx_test_projects/filterbank_ip
    --  set_property -dict [list CONFIG.Component_Name {PSSFBReorderMem} CONFIG.Memory_Type {Simple_Dual_Port_RAM} CONFIG.Assume_Synchronous_Clk {true} CONFIG.Write_Width_A {192} CONFIG.Write_Depth_A {128} CONFIG.Read_Width_A {192} CONFIG.Operating_Mode_A {NO_CHANGE} CONFIG.Enable_A {Always_Enabled} CONFIG.Write_Width_B {192} CONFIG.Read_Width_B {192} CONFIG.Operating_Mode_B {READ_FIRST} CONFIG.Enable_B {Always_Enabled} CONFIG.Register_PortA_Output_of_Memory_Primitives {false} CONFIG.Register_PortB_Output_of_Memory_Primitives {true} CONFIG.Fill_Remaining_Memory_Locations {true} CONFIG.Port_B_Clock {100} CONFIG.Port_B_Enable_Rate {100} CONFIG.Collision_Warnings {GENERATE_X_ONLY} CONFIG.Disable_Collision_Warnings {true} CONFIG.Disable_Out_of_Range_Warnings {true}] [get_ips PSSFBReorderMem]
    component PSSFBReorderMem
    port (
        clka  : in std_logic;
        wea   : in std_logic_vector(0 downto 0);
        addra : in std_logic_vector(6 downto 0);
        dina  : in std_logic_vector(191 downto 0);
        clkb  : in std_logic;
        addrb : in std_logic_vector(6 downto 0);
        doutb : out std_logic_vector(191 downto 0));
    end component;
    
    signal wrData96 : std_logic_vector(95 downto 0);
    signal FBmemRdData : t_slv_96_arr(11 downto 0);
    signal FBmemFIRTaps : t_slv_18_arr(11 downto 0);
    
    -- The first index in fbtype is for the number of filters = 12 (6 channels * 2[real+imaginary]).
    -- The second index is for the number of FIR taps.
    type fbtype is array(11 downto 0) of t_slv_8_arr(11 downto 0); 
    signal FBRdData : fbtype;
    signal FIRDout : t_slv_16_arr(11 downto 0);
    signal fftIndex : t_slv_6_arr(5 downto 0);
    
    signal fftRealOut : t_slv_16_arr(5 downto 0);
    signal fftImagOut : t_slv_16_arr(5 downto 0);
    signal fftvalidOut : std_logic_vector(5 downto 0) := "000000";
    
    signal startAdv : std_logic_vector(31 downto 0);
    signal validDel1, validDel2 : std_logic := '0';
    signal startFFT : std_logic := '0';
    
    signal reorderDout : std_logic_vector(191 downto 0);
    signal reorderWE : std_logic_vector(0 downto 0);
    signal reorderWrAddr : std_logic_vector(5 downto 0);
    signal reorderWrAddrFull : std_logic_vector(6 downto 0);
    signal reorderRdAddr : std_logic_vector(5 downto 0);
    signal reorderRdAddrFull : std_logic_vector(6 downto 0);
    signal bufSelectWr, bufSelectRd : std_logic := '0';
    signal reorderDin : std_logic_vector(191 downto 0);
    signal rdRunning : std_logic := '0';
    signal rdRunningDel2, rdRunningDel1 : std_logic := '0';
    signal validOutDel1 : std_logic := '0';
    signal bufSelectRdDel1, bufSelectRdDel2 : std_logic := '0';
    
begin
    
    ------------------------------------------------------------------------------------
    -- 1. Input Memory
    -- ---------------
    
    wrData96 <= data5_i(1) & data5_i(0) & data4_i(1) & data4_i(0) & data3_i(1) & data3_i(0) & data2_i(1) & data2_i(0) & data1_i(1) & data1_i(0) & data0_i(1) & data0_i(0);

    cmem : entity filterbanks_lib.PSSFBMem
    generic map (
        TAPS => 12)  -- Note only partially parameterized; modification needed to support anything other than 12.
    port map (
        clk         => clk,
        FIRTapUse_i => FIRTapUse_i,   -- in std_logic; FIR Taps are double buffered, choose which set of TAPs to use.
        -- Write data for the start of the chain
        wrData_i    => wrData96,      -- in(95:0);
        wrEn_i      => valid_i,       -- in std_logic; should be a burst of 4096 clocks.
        -- Read data, comes out 2 clocks after the first write.
        rd_data_o   => FBmemRdData,   -- out array96bit_type(TAPS-1 downto 0); -- 64 bits wide, 12 taps simultaneously; First sample is wr_data_i delayed by 1 clock. 
        coef_o      => FBmemFIRTaps,  -- out array18bit_type(TAPS-1 downto 0); -- 18 bits per filter tap.
        -- Writing FIR Taps
        FIRTapData_i   => FIRTapData_i,   -- in(17:0);  -- For register writes of the filtertaps.
        FIRTapData_o   => FIRTapData_o,   -- out(17:0); -- For register reads of the filtertaps. 3 cycle latency from FIRTapAddr_i
        FIRTapAddr_i   => FIRTapAddr_i,   -- in(11:0);  -- 64 * 12 filter taps = 768 total.
        FIRTapWE_i     => FIRTapWE_i,     -- in std_logic;
        FIRTapClk      => FIRTapClk,      -- in std_logic;
        FIRTapSelect_i => FIRTapSelect_i  -- in std_logic; FIR Taps are double buffered; this selects the buffer to access for registers. Choose which buffer to use with FIRTapUse_i
    );
    
    -------------------------------------------------------------------------------------
    -- 2. FIR filter
    -- -------------
    -- 12 instances, 6 channels * (real + imaginary). Same filter taps used for all.
    -- PISA low.CBF processes simultaneously 2 (real+imaginary) * 3 (stations) * 2 (polarisations) = 12
    -- 
    
    CsampleGen : for j in 0 to 11 generate  -- 12 filters
        coefGen : for k in 0 to 11 generate  -- 12 taps
            FBRdData(j)(k) <= FBmemRdData(k)((j*8 + 7) downto (j*8));
        end generate;
    end generate;
    
    sampleGen : for j in 0 to 11 generate
            
        FIR : entity filterbanks_lib.fb_DSP
        generic map (
            TAPS => 12)  -- The module instantiates this number of DSPs
        port map (
            clk    => clk,
            data_i => FBRdData(j),  -- in array8bit_type(11 downto 0);
            coef_i => FBmemFIRTaps, -- in array18bit_type(11 downto 0);
            data_o => FIRDout(j)    -- out(15:0)
        );
    
    end generate;
    
    -------------------------------------------------------------------------------------
    -- 3. FFT
    -- -----------------
    -- 6 x 64 point FFTs.
    
    process(clk)
    begin
        if rising_edge(clk) then
            validDel1 <= valid_i;
            validDel2 <= validDel1;
            if validDel1 = '1' and validDel2 = '0' then
                startAdv(0) <= '1';
            else
                startAdv(0) <= '0';
            end if;
            
            startAdv(31 downto 1) <= startAdv(30 downto 0);
            startFFT <= startAdv(12); -- Delay accounts for the delay through the FIR filter 
            
        end if;
    end process;
    
    
    fftgen : for j in 0 to 5 generate
        
        fft64 : entity filterbanks_lib.PSSFFTwrapper
        port map (
            clk  => clk,
            -- Input
            real_i  => FIRDout(j*2),     -- in(15:0); 16 bit real data
            imag_i  => FIRDout(j*2 + 1), -- in(15:0); 16 bit imaginary data
            start_i => startFFT,         -- in std_logic; pulse high; one clock in advance of the data 
            -- Output
            real_o  => fftRealOut(j), -- out(15:0);
            imag_o  => fftImagOut(j), -- out(15:0);
            index_o => fftIndex(j),   -- out(5:0);
            valid_o => fftvalidOut(j) -- out std_logic
        );
    
    end generate;
    
    -------------------------------------------------------------------------------------
    -- 4. Reorder the output from bit-reversed to the central 54 channels, low to high frequency.
    -- Uses a simple dual port BRAM double buffer.
      
    process(clk)
    begin
        if rising_edge(clk) then
        
            if (fftvalidOut(0) = '1' and (signed(fftIndex(0)) > -28) and (signed(fftIndex(0)) < 27)) then
                reorderWE(0) <= '1';
            else
                reorderWE(0) <= '0';
            end if;
            reorderWrAddr <= std_logic_vector(signed(fftIndex(0)) + 27);
            reorderDin <= fftImagOut(5) & fftRealOut(5) & fftImagOut(4) & fftRealOut(4) & fftImagOut(3) & fftRealOut(3) & fftImagOut(2) & fftRealOut(2) & fftImagOut(1) & fftRealOut(1) & fftImagOut(0) & fftRealOut(0);
            
            -- Falling edge of validOut triggers reading of the data from the memory
            validOutDel1 <= fftvalidOut(0);
            if fftvalidOut(0) = '0' and validOutDel1 = '1' then
                reorderRdAddr <= "000000";
                bufSelectWr <= not bufSelectWr;
                bufSelectRd <= bufSelectWr;
                rdRunning <= '1';
            elsif rdRunning = '1' then
                reorderRdAddr <= std_logic_vector(unsigned(reorderRdAddr) + 1);
                -- read address runs from 0 to 53
                if unsigned(reorderRdAddr) = 53 then
                   rdRunning <= '0';
                end if;
            end if;
            rdRunningDel1 <= rdRunning;
            rdRunningDel2 <= rdRunningDel1;
            bufSelectRdDel1 <= bufSelectRd;
            bufSelectRdDel2 <= bufSelectRdDel1;
        end if;
    end process;
    
    reorderWrAddrFull <= bufSelectWr & reorderWrAddr;
    reorderRdAddrFull <= bufSelectRd & reorderRdAddr;
    
    reorderRAM : PSSFBReorderMem
    port map (
        clka  => clk,
        wea   => reorderWE,         -- in std_logic_vector(0 downto 0);
        addra => reorderWrAddrFull, -- in(6:0);
        dina  => reorderDin,        -- in(95:0);
        clkb  => clk,
        addrb => reorderRdAddrFull, -- in(6:0);
        doutb => reorderDout        -- out(95:0)
    );

    process(clk)
    begin
        if rising_edge(clk) then
            data0_o(0) <= reorderDout(15 downto 0);
            data0_o(1) <= reorderDout(31 downto 16);
            data1_o(0) <= reorderDout(47 downto 32);
            data1_o(1) <= reorderDout(63 downto 48);
            data2_o(0) <= reorderDout(79 downto 64);
            data2_o(1) <= reorderDout(95 downto 80);
            data3_o(0) <= reorderDout(111 downto 96);
            data3_o(1) <= reorderDout(127 downto 112);
            data4_o(0) <= reorderDout(143 downto 128);
            data4_o(1) <= reorderDout(159 downto 144);
            data5_o(0) <= reorderDout(175 downto 160);
            data5_o(1) <= reorderDout(191 downto 176);
            valid_o <= rdRunningDel2;
        end if;
    end process;    
    
end Behavioral;
