-------------------------------------------------------------------------------
-- Title      : Mid Term Accumulator Registers
-- Project    : 
-------------------------------------------------------------------------------
-- File       : mta_regs_pkg.vhd
-- Author     : William Kamp  <william.kamp@aut.ac.nz>
-- Company    : High Performance Computing Research Lab, Auckland University of Technology
-- Created    : 2018-01-05
-- Last update: 2018-01-08
-- Platform   : 
-- Standard   : VHDL'08
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Copyright (c) 2018 High Performance Computing Research Lab, Auckland University of Technology
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2018-01-05  1.0      will    Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;

package mta_regs_pkg is

    type t_cci_ram_wr_reg is record
        clk        : std_logic;
        reset      : std_logic;
        address    : unsigned(31 downto 0);
        wr_req     : std_logic;
        cci_factor : std_logic_vector(31 downto 0);
    end record t_cci_ram_wr_reg;

    -- autogen start decl
 --------------------------------------------------
 -- Auto-generated code below. You should not edit.
 -- Generated Mon Jan  8 15:10:19 2018
 --------------------------------------------------
type t_cci_ram_wr_reg_a is array(natural range <>) of t_cci_ram_wr_reg;

constant T_CCI_RAM_WR_REG_ZERO : t_cci_ram_wr_reg := (
	clk => '0',
	reset => '0',
	address => (others => '0'),
	wr_req => '0',
	cci_factor => (others => '0')
	);

constant T_CCI_RAM_WR_REG_DONT_CARE : t_cci_ram_wr_reg := (
	clk => '-',
	reset => '-',
	address => (others => '-'),
	wr_req => '-',
	cci_factor => (others => '-')
	);

constant T_CCI_RAM_WR_REG_SLV_WIDTH : natural := 67;

subtype t_cci_ram_wr_reg_slv is std_logic_vector(66 downto 0);
function to_slv (rec : t_cci_ram_wr_reg) return t_cci_ram_wr_reg_slv;

function from_slv (slv : std_logic_vector) return t_cci_ram_wr_reg;

 ------------------------------------------------------
 -- End of Autogenerated code. You may add yours below.
 ------------------------------------------------------
    -- autogen end decl

end package mta_regs_pkg;

package body mta_regs_pkg is

    -- autogen start body
 --------------------------------------------------
 -- Auto-generated code below. You should not edit.
 -- Generated Mon Jan  8 15:10:19 2018
 --------------------------------------------------
function to_slv (rec : t_cci_ram_wr_reg) return t_cci_ram_wr_reg_slv is
    variable slv : std_logic_vector(66 downto 0);
begin
    slv(31 downto 0) := rec.cci_factor;
    slv(32) := rec.wr_req;
    slv(64 downto 33) := std_logic_vector(rec.address);
    slv(65) := rec.reset;
    slv(66) := rec.clk;
return slv;
end function to_slv;

function from_slv (slv : std_logic_vector) return t_cci_ram_wr_reg is
    variable rec : t_cci_ram_wr_reg;
begin
    rec.cci_factor := slv(31 downto 0);
    rec.wr_req := slv(32);
    rec.address := unsigned(slv(64 downto 33));
    rec.reset := slv(65);
    rec.clk := slv(66);
return rec;
end function from_slv;

 ------------------------------------------------------
 -- End of Autogenerated code. You may add yours below.
 ------------------------------------------------------
    -- autogen end body

end package body mta_regs_pkg;
