-------------------------------------------------------------------------------
--
-- Copyright (C) 2017
-- CSIRO
--
-- This program is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
--
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with this program.  If not, see <http://www.gnu.org/licenses/>.
--
-------------------------------------------------------------------------------

-- Purpose: <fpga_name>_bus_top specific constants and functions
--
-- Description:
--
-- Remarks:
--  This file was automatically generated by ARGS from <fpga_name>.peripheral.yaml

LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;

PACKAGE <fpga_name>_bus_pkg IS

    CONSTANT c_nof_lite_slaves  : NATURAL := <nof_lite_slaves>;
    CONSTANT c_nof_full_slaves  : NATURAL := <nof_full_slaves>;

    CONSTANT c_data_w   : NATURAL := 32;
    CONSTANT c_addr_w   : NATURAL := 32;
    CONSTANT c_strb_w   : NATURAL := 4;

    -- Lite slave port indexes
<{LITE}>    CONSTANT c_{}_lite_index<tabs>: NATURAL := {};

    -- Full slave port indexes
<{FULL}>    CONSTANT c_{}_full_index<tabs>: NATURAL := {};

END <fpga_name>_bus_pkg;

PACKAGE BODY <fpga_name>_bus_pkg IS

END <fpga_name>_bus_pkg;