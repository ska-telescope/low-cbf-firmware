----------------------------------------------------------------------------------
-- Company: CSIRO 
-- Engineer: David Humphrey (dave.humphrey@csiro.au)
-- 
-- Create Date: 18.07.2019
-- Module Name: IC_outputMux - Behavioral
-- 
-- Description 
-- -----------
--   + Watches for notifications of packets that are available, and puts them into a FIFO
--   + Requests transmission of packets from the input modules, and muxes the data and valid signal onto the output bus.
--
-- Details
-- -------
--   Notifications are generated by all the input buffers. In the IC_top module, they are muxed down
--  to a single bus which goes to all the output buffers.
--  Notifications contain 
--   * The destination address for the packet (i_NotificationAddress). The address includes the XYZ coordinates of the destination FPGA,
--     as well as the signal chain port it is going to.
--   * The location in the input buffer memory (the "block") where the packet starts (i_NotificationBlock)
--   * The input port that the notification came from (i_NotificationPort)
--  This module looks at the destination address and compares with the destination address and port configured for this output mux.
--  If it matches this module, then the notification goes into the notification FIFO.
--  The FIFO stores the input port and the block.
--  The last four entries in the FIFO are stored in registers so that they can be read out of order.
--  This means that if an input port is busy sending a packet somewhere else, then we can request a packet from a different input
--  port.
--  The valid output from all the input ports is visible in this module, so we can detect if an input port is busy sending data to
--  some other output port.
--  When we need more data, the block and input port are placed on the request bus. 
--  After placing the data on the request bus, we watch that input port (i_packetDest(port)) for our address, and if it
--  matches, we forward the data from that port.
--  If it doesn't match, then the input port must have allocated itself to another output port. In this case, this module withdraws 
--  its request and can request from another input port (if there are other packets waiting to be sent).
--  Note : The input side ports should enforce a minimum packet length of 8 words, to avoid allocating to an output port
--  that has dropped the request.
--
-- "PORTSUSED"
-- -------
--  The generic PORTSUSED allows for ports to be masked out of the output multiplexer in order to save resources.
--  If an input port that is masked out makes a request to this output port, then the o_inputPortInvalid flag is raised.
--
-- Addressing
-- ----------
-- The first (64 bit) word of each packet must contain :
--
--   DEST    SRC1     SRC2    SRC3     PacketTYPE
-- (63:52)  (51:40)  (39:28) (27:16)  (15:8)
-- 
-- Each address (DEST, SRC1, SRC2, SRC3) is made up of 
--  (11:8) = Y coordinate
--  (7:4) = X coordinate
--  (3:0) = Z coordinate
--
-- Packets travel through FPGAs in in the order : SRC3 -> SRC2 -> SRC1 -> DEST
-- If there are less than 3 hops to the destination, then the unused addresses are 0xfff
-- e.g. a single hop packet would have SRC3 = SRC2 = 0xfff
-- 
-- The interconnect module has output ports which go to each possible destination. 
-- The output ports are numbered as :
--  0-7 : Z connect (e.g. port 3 sends data over the fiber going to the FPGA with Z = 3 and the same X,Y coordinates as this FPGA)
--  8-13 : X connect
--  14-19 : Y connect
--  20 up : The signal processing chain in this FPGA, identified as (20 + packetType)
-- 
-- Why allow out-of-order reads ?
-- ------------------------------
-- This is to ensure the optical links are used efficiently, since the destination port for a given
-- packet could be busy with a packet from another source port, temporarily blocking this port. 
-- Blocking is statistically likely to occur for a non-negligible portion of the time, impacting the 
-- overall performance of the interconnect, since the average rate into the URAM cannot exceed the average rate out without
-- causing packets to be lost. By allowing packets other than the oldest packet in the buffer to be read when the destination
-- port is ready, the probability of blocking is significantly reduced.
--  
----------------------------------------------------------------------------------

library common_lib;
use common_lib.common_pkg.all;
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
Library xpm;
use xpm.vcomponents.all;

entity IC_outputMux is
    generic(
        -- 0 = 3 FPGAs (X x Y x Z = 1x1x3), 1 = 12 FPGAs (X x Y x Z = 1x6x2), 2 = etc....
        -- See confluence page (perentie -> Model development -> packetised model overview -> model configuration)    
        ARRAYRELEASE : integer range 0 to 5 := 0;
        -- PortsUsed allows input side ports to be masked out from the multiplexer to save resources. 
        -- Set bits to 0 to mask a port.
        PORTSUSED : std_logic_vector(31 downto 0) := x"ffffffff";
        OUTPUTMUX : std_logic_vector(4 downto 0);  -- index of this output mux
        FIBEROUTPUT : std_logic := '1';  -- this module sends data to a GTY
        DROPADDRWORD : std_logic := '0'  -- drop the first word of the packet (the address word). Signal chain modules don't expect the address word.
    );
    port(
        -- Everything is on a single clock (about 400 MHz)
        i_IC_clk : in std_logic;
        i_rst : in std_logic;
        -- Configuration information
        i_myAddr : in std_logic_vector(11 downto 0);   -- X,Y and Z coordinates of this FPGA in the array, used for routing.
        i_destAddr : in std_logic_vector(11 downto 0); -- X,Y and Z coordinates of the place this output mux sends data to.
        i_destPort : in std_logic_vector(3 downto 0);  -- signal chain port this output mux sends data to. Only used if i_myAddr = i_destAddr, (i.e. when packets coming to this mux are destined for this FPGA).
        -- Packet Data being streamed out by the input side modules 
        i_packetData  : in t_slv_64_arr(31 downto 0);      -- 
        i_packetOutputMux : in t_slv_5_arr(31 downto 0);   -- Destination output MUX for this packet (i.e. send the packet through this module if i_packetOutputMux = OUTPUTMUX).
        i_packetValid : in std_logic_vector(31 downto 0);
        -- Notification from input ports of packets being available at a particular block in a buffer 
        -- These go to a FIFO in this module, if the destination address matches i_destAddr, i_destPort.
        i_NotificationAddress : in std_logic_vector(15 downto 0); -- destination address for this packet, (11:0) = XYZ coordinates, (15:12) = signal chain port. 
        i_NotificationBlock   : in std_logic_vector(4 downto 0);  -- the block in the buffer that the packet is stored at.
        i_NotificationPort    : in std_logic_vector(4 downto 0);  -- the input port that this notification comes from.
        i_NotificationValid   : in std_logic;
        -- Requests out to the input ports
        o_RequestBlock : out std_logic_vector(4 downto 0); -- Block in the buffer that we want to get data from.
        o_RequestPort  : out std_logic_vector(4 downto 0); -- The input port that data is being requested from
        o_RequestValid : out std_logic;                    -- o_block and o_port are valid. 
        -- The packets
        o_data  : out std_logic_vector(63 downto 0);
        o_sop   : out std_logic;
        o_valid : out std_logic;
        -- Status
        i_clrErrorCounts : in std_logic;
        o_errCounts : out std_logic_vector(7 downto 0)  -- (3:0) = fifo full, bit(3) is sticky; (7:4) = input port invalid count, bit(7) is sticky.
    );
end IC_outputMux;

architecture Behavioral of IC_outputMux is

    type rd_fsm_type is (idle, getAvailable, waitRequest, sendData);
    signal rd_fsm, rd_fsm_del : rd_fsm_type := idle;

    -- 4 entry fifo built from registers so we can read any entry when we need to
    signal fifoRd : std_logic;
    signal fifoRdEntry : std_logic_vector(1 downto 0);
    signal fifoUsed, fifoUsedRdfsm : std_logic_vector(3 downto 0);
    signal fifoEntry0, fifoEntry1, fifoEntry2, fifoEntry3 : std_logic_vector(9 downto 0);
    signal fifoCompact : std_logic;
    -- 4 entry fifo is fed from "mainFifo", which is 32 deep.
    signal mainFifoRdData : std_logic_vector(9 downto 0);
    signal mainFifoRdEn : std_logic := '0';
    signal mainFifoEmpty : std_logic;
    
    COMPONENT IC_omux_FIFO
    PORT (
        clk   : IN STD_LOGIC;
        srst  : IN STD_LOGIC;
        din   : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
        wr_en : IN STD_LOGIC;
        rd_en : IN STD_LOGIC;
        dout  : OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
        full  : OUT STD_LOGIC;
        empty : OUT STD_LOGIC;
        wr_rst_busy : OUT STD_LOGIC;
        rd_rst_busy : OUT STD_LOGIC);
    END COMPONENT;

    signal selectedPacketData : std_logic_vector(63 downto 0);
    signal maskedPacketData : t_slv_64_arr(31 downto 0);
    signal selectedOutputMux : std_logic_vector(4 downto 0);
    signal selectedPacketValid : std_logic;
    signal validSel0, validSel1, validSel2, validSel3 : std_logic;
    signal requestPort : std_logic_vector(4 downto 0);
    signal mainFifoDin : std_logic_vector(9 downto 0);
    signal mainFifoWrEn : std_logic;
    signal mainFifoFull : std_logic;
    signal wr_rst_busy, rd_rst_busy : std_logic;
    signal selectedPortPossible : std_logic;
    signal oinputPortInvalid : std_logic;
    signal ostatFifoFull : std_logic;
    signal anyPortInvalid : std_logic := '0';
    signal portInvalidCount : std_logic_vector(2 downto 0) := "000";
    signal anyfifoFull : std_logic := '0';
    signal fifoFullCount : std_logic_vector(2 downto 0) := "000";
    signal validDel : std_logic;
    signal selectedPacketValidDel : std_logic := '0';
    signal valid_int : std_logic;
    
begin
    
    ------------------------------------------------------------------------------------------------
    -- Fifo for notifications
    ------------------------------------------------------------------------------------------------
    
    process(i_IC_clk)
    begin
        if rising_edge(i_IC_clk) then
            
            -- Four entry shift register for the output of the notification fifo, so we can choose 
            -- any of up to four packets which are available from the input ports.
            --
            -- The shift register is built out of 
            --
            if i_rst = '1' then
                fifoUsed <= "0000";
                mainFifoRdEn <= '0';
            elsif fifoRd = '1' then
                if fifoRdEntry = "00" then
                    fifoUsed(0) <= '0';
                elsif fifoRdEntry = "01" then
                    fifoUsed(1) <= '0';
                elsif fifoRdEntry = "10" then
                    fifoUsed(2) <= '0';
                else
                    fifoUsed(3) <= '0';
                end if;
                if mainFifoRdEn = '1' then
                    mainFifoRdEn <= '0';
                    if fifoUsed = "0000" then
                        fifoEntry0 <= mainFifoRdData;
                        fifoUsed(0) <= '1';
                    elsif fifoUsed(3 downto 1) = "000" then
                        fifoEntry1 <= mainFifoRdData;
                        fifoUsed(1) <= '1';
                    elsif fifoUsed(3 downto 2) = "00" then
                        fifoEntry2 <= mainFifoRdData;
                        fifoUsed(2) <= '1';
                    else
                        fifoEntry3 <= mainFifoRdData;
                        fifoUsed(3) <= '1';
                    end if;
                end if;
            elsif mainFifoRdEn = '1' then
                mainFifoRdEn <= '0';
                if fifoUsed = "0000" then
                    fifoEntry0 <= mainFifoRdData;
                    fifoUsed(0) <= '1';
                elsif fifoUsed(3 downto 1) = "000" then
                    fifoEntry1 <= mainFifoRdData;
                    fifoUsed(1) <= '1';
                elsif fifoUsed(3 downto 2) = "00" then
                    fifoEntry2 <= mainFifoRdData;
                    fifoUsed(2) <= '1';
                else
                    fifoEntry3 <= mainFifoRdData;
                    fifoUsed(3) <= '1';
                end if;
            elsif fifoCompact = '0' and fifoUsed /= "0000" then
                mainFifoRdEn <= '0';
                if fifoUsed(0) = '0' and fifoUsed(3 downto 1) /= "000" then
                    fifoEntry0 <= fifoEntry1;
                    fifoEntry1 <= fifoEntry2;
                    fifoEntry2 <= fifoEntry3;
                    fifoUsed(3 downto 0) <= '0' & fifoUsed(3 downto 1);
                elsif fifoUsed(1) = '0' and fifoUsed(3 downto 2) /= "00" then
                    fifoEntry1 <= fifoEntry2;
                    fifoEntry2 <= fifoEntry3;
                    fifoUsed(3 downto 1) <= '0' & fifoUsed(3 downto 2);
                elsif fifoUsed(2) = '0' and fifoUsed(3) /= '0' then
                    fifoEntry2 <= fifoEntry3;
                    fifoUsed(3 downto 2) <= '0' & fifoUsed(3);
                end if;
            elsif fifoUsed(3) = '0' and mainFifoEmpty = '0' and mainFifoRdEn = '0' then
                mainFifoRdEn <= '1';
            end if;
            
            -- Write notifications to the mainFifo if
            --     - The destination address is the address of this FPGA (i_myAddr) and the destination signal chain port is the port his mux is connected to (i_destPort)
            --  or - The destination address is the address this mux is sending to (i_destAddr) and this mux is sending to a fiber output (i.e. not to a signal chain output)
            if (((i_NotificationAddress(11 downto 0) = i_myAddr and i_NotificationAddress(15 downto 12) = i_destPort) or 
                (i_NotificationAddress(11 downto 0) = i_destAddr and (FIBEROUTPUT = '1'))) and i_NotificationValid = '1') then
                mainFifoWrEn <= '1';
            else
                mainFifoWrEn <= '0';
            end if;
            mainFifoDin <= i_notificationPort & i_notificationBlock;
            ostatFifoFull <= mainFifoFull;
            
        end if;
    end process;
    
    
    -- Only read from the fifo is the output is compacted.
    -- Otherwise we could read but have the location of the entry we are reading move.
    fifoCompact <= '1' when fifoUsed = "0001" or fifoUsed = "0011" or fifoUsed = "0111" or fifoUsed = "1111" else '0';
    
    xpm_fifo_sync_inst : xpm_fifo_sync
    generic map (
        DOUT_RESET_VALUE => "0",    -- String, Reset value of read data path.
        ECC_MODE => "no_ecc",       -- String, Allowed values: no_ecc, en_ecc.
        FIFO_MEMORY_TYPE => "distributed", -- String, Allowed values: auto, block, distributed. 
        FIFO_READ_LATENCY => 0,     -- Integer, Range: 0 - 10. Must be 0 for first READ_MODE = "fwft" (first word fall through).    
        FIFO_WRITE_DEPTH => 32,     -- Integer, Range: 16 - 4194304. Defines the FIFO Write Depth. Must be power of two.
        FULL_RESET_VALUE => 0,      -- Integer, Range: 0 - 1. Sets full, almost_full and prog_full to FULL_RESET_VALUE during reset
        PROG_EMPTY_THRESH => 10,    -- Integer, Range: 3 - 4194301.Specifies the minimum number of read words in the FIFO at or below which prog_empty is asserted.
        PROG_FULL_THRESH => 10,     -- Integer, Range: 5 - 4194301. Specifies the maximum number of write words in the FIFO at or above which prog_full is asserted.
        RD_DATA_COUNT_WIDTH => 1,   -- Integer, Range: 1 - 23. Specifies the width of rd_data_count. To reflect the correct value, the width should be log2(FIFO_READ_DEPTH)+1. FIFO_READ_DEPTH = FIFO_WRITE_DEPTH*WRITE_DATA_WIDTH/READ_DATA_WIDTH         
        READ_DATA_WIDTH => 10,      -- Integer, Range: 1 - 4096. Defines the width of the read data port, dout
        READ_MODE => "fwft",        -- String, Allowed values: std, fwft. Default value = std.
        --SIM_ASSERT_CHK => 0,        -- DECIMAL; 0=disable simulation messages, 1=enable simulation messages
        USE_ADV_FEATURES => "0000", -- String
        -- |---------------------------------------------------------------------------------------------------------------------|
        -- | Enables data_valid, almost_empty, rd_data_count, prog_empty, underflow, wr_ack, almost_full, wr_data_count,         |
        -- | prog_full, overflow features.                                                                                       |
        -- |                                                                                                                     |
        -- |   Setting USE_ADV_FEATURES[0] to 1 enables overflow flag;     Default value of this bit is 1                        |
        -- |   Setting USE_ADV_FEATURES[1]  to 1 enables prog_full flag;    Default value of this bit is 1                       |
        -- |   Setting USE_ADV_FEATURES[2]  to 1 enables wr_data_count;     Default value of this bit is 1                       |
        -- |   Setting USE_ADV_FEATURES[3]  to 1 enables almost_full flag;  Default value of this bit is 0                       |
        -- |   Setting USE_ADV_FEATURES[4]  to 1 enables wr_ack flag;       Default value of this bit is 0                       |
        -- |   Setting USE_ADV_FEATURES[8]  to 1 enables underflow flag;    Default value of this bit is 1                       |
        -- |   Setting USE_ADV_FEATURES[9]  to 1 enables prog_empty flag;   Default value of this bit is 1                       |
        -- |   Setting USE_ADV_FEATURES[10] to 1 enables rd_data_count;     Default value of this bit is 1                       |
        -- |   Setting USE_ADV_FEATURES[11] to 1 enables almost_empty flag; Default value of this bit is 0                       |
        -- |   Setting USE_ADV_FEATURES[12] to 1 enables data_valid flag;   Default value of this bit is 0                       |
        WAKEUP_TIME => 0,          -- Integer, Range: 0 - 2. 0 = Disable sleep 
        WRITE_DATA_WIDTH => 10,    -- Integer, Range: 1 - 4096. Defines the width of the write data port, din             
        WR_DATA_COUNT_WIDTH => 1   -- Integer, Range: 1 - 23. Specifies the width of wr_data_count. To reflect the correct value, the width should be log2(FIFO_WRITE_DEPTH)+1.   |
    )
    port map (
        almost_empty => open, -- 1-bit output: Almost Empty : When asserted, this signal indicates that only one more read can be performed before the FIFO goes to empty.
        almost_full => open,  -- 1-bit output: Almost Full: When asserted, this signal indicates that only one more write can be performed before the FIFO is full.
        data_valid => open,   -- 1-bit output: Read Data Valid: When asserted, this signal indicates that valid data is available on the output bus (dout).
        dbiterr => open,      -- 1-bit output: Double Bit Error: Indicates that the ECC decoder detected a double-bit error and data in the FIFO core is corrupted.
        dout => mainFifoRdData,  -- READ_DATA_WIDTH-bit output: Read Data: The output data bus is driven when reading the FIFO.
        empty => mainFifoEmpty,  -- 1-bit output: Empty Flag: When asserted, this signal indicates that
                                 -- the FIFO is empty. Read requests are ignored when the FIFO is empty, initiating a read while empty is not destructive to the FIFO.
        full => mainFifofull,    -- 1-bit output: Full Flag: When asserted, this signal indicates that the FIFO is full. Write requests are ignored when the FIFO is full,
                                 -- initiating a write when the FIFO is full is not destructive to the contents of the FIFO.
        overflow => open,   -- 1-bit output: Overflow: This signal indicates that a write request (wren) during the prior clock cycle was rejected, because the FIFO is
                            -- full. Overflowing the FIFO is not destructive to the contents of the FIFO.
        prog_empty => open, -- 1-bit output: Programmable Empty: This signal is asserted when the number of words in the FIFO is less than or equal to the programmable
                            -- empty threshold value. It is de-asserted when the number of words in the FIFO exceeds the programmable empty threshold value.
        prog_full => open,  -- 1-bit output: Programmable Full: This signal is asserted when the number of words in the FIFO is greater than or equal to the
                            -- programmable full threshold value. It is de-asserted when the number of words in the FIFO is less than the programmable full threshold value.
        rd_data_count => open,      -- RD_DATA_COUNT_WIDTH-bit output: Read Data Count: This bus indicates the number of words read from the FIFO.
        rd_rst_busy => rd_rst_busy, -- 1-bit output: Read Reset Busy: Active-High indicator that the FIFO read domain is currently in a reset state.
        sbiterr => open,            -- 1-bit output: Single Bit Error: Indicates that the ECC decoder detected and fixed a single-bit error.
        underflow => open,          -- 1-bit output: Underflow: Indicates that the read request (rd_en) during the previous clock cycle was rejected because the FIFO is empty. Under flowing the FIFO is not destructive to the FIFO.
        wr_ack => open,             -- 1-bit output: Write Acknowledge: This signal indicates that a write request (wr_en) during the prior clock cycle is succeeded.
        wr_data_count => open,      -- WR_DATA_COUNT_WIDTH-bit output: Write Data Count: This bus indicates the number of words written into the FIFO.
        wr_rst_busy => wr_rst_busy, -- 1-bit output: Write Reset Busy: Active-High indicator that the FIFO write domain is currently in a reset state.
        din => mainFifoDin,         -- WRITE_DATA_WIDTH-bit input: Write Data: The input data bus used when writing the FIFO.
        injectdbiterr => '0',       -- 1-bit input: Double Bit Error Injection: Injects a double bit error if the ECC feature is used on block RAMs or UltraRAM macros.
        injectsbiterr => '0',       -- 1-bit input: Single Bit Error Injection: Injects a single bit error if the ECC feature is used on block RAMs or UltraRAM macros.
        rd_en => mainFifoRdEn,      -- 1-bit input: Read Enable: If the FIFO is not empty, asserting this signal causes data (on dout) to be read from the FIFO. Must be held active-low when rd_rst_busy is active high.
        rst => i_rst,               -- 1-bit input: Reset.
        sleep => '0',               -- 1-bit input: Dynamic power saving: If sleep is High, the memory/fifo block is in power saving mode.
        wr_clk => i_IC_clk,         -- 1-bit input: Write clock: Used for write operation. wr_clk must be a free running clock.
        wr_en => mainFifoWrEn       -- bit input: Write Enable: If the FIFO is not full, asserting this signal causes data (on din) to be written to the FIFO. Must be held active-low when rst or wr_rst_busy is active high.
    );
    
    --------------------------------------------------------------------------------------------------
    -- Read the notification FIFO, generate requests to the input ports, 
    -- and mux the output data onto o_valid, o_data.
    
    process(i_IC_clk)
        variable sel0, sel1, sel2, sel3 : std_logic_vector(4 downto 0);
    begin
        if rising_edge(i_IC_clk) then
            case rd_fsm is
                when idle =>
                    if fifoCompact = '1' then
                        rd_fsm <= getAvailable;
                    end if;
                    fifoUsedRdfsm <= fifoUsed;
                    sel0 := fifoEntry0(9 downto 5);
                    sel1 := fifoEntry1(9 downto 5);
                    sel2 := fifoEntry2(9 downto 5);
                    sel3 := fifoEntry3(9 downto 5);
                    validSel0 <= i_PacketValid(to_integer(unsigned(sel0)));
                    validSel1 <= i_PacketValid(to_integer(unsigned(sel1)));
                    validSel2 <= i_PacketValid(to_integer(unsigned(sel2)));
                    validSel3 <= i_PacketValid(to_integer(unsigned(sel3)));
                    o_RequestValid <= '0'; 
                    o_RequestBlock <= "00000";
                    RequestPort <= "00000";
                    fifoRdEntry <= "00";
                    
                when getAvailable =>
                    if fifoUsedRdfsm(0) = '1' and validSel0 = '0' then -- Get data from input buffer sel0 
                        rd_fsm <= waitRequest;
                        o_RequestBlock <= fifoEntry0(4 downto 0);
                        RequestPort <= fifoEntry0(9 downto 5);
                        fifoRdEntry <= "00";
                        o_RequestValid <= '1';
                    elsif fifoUsedRdfsm(1) = '1' and validSel1 = '0' then 
                        rd_fsm <= waitRequest;
                        o_RequestBlock <= fifoEntry1(4 downto 0);
                        RequestPort <= fifoEntry1(9 downto 5);
                        fifoRdEntry <= "01";
                        o_RequestValid <= '1';
                    elsif fifoUsedRdfsm(2) = '1' and validSel2 = '0' then
                        rd_fsm <= waitRequest;
                        o_RequestBlock <= fifoEntry2(4 downto 0);
                        RequestPort <= fifoEntry2(9 downto 5);
                        fifoRdEntry <= "10";
                        o_RequestValid <= '1';
                    elsif fifoUsedRdfsm(3) = '1' and validSel3 = '0' then
                        rd_fsm <= waitRequest;
                        o_RequestBlock <= fifoEntry3(4 downto 0);
                        RequestPort <= fifoEntry3(9 downto 5);
                        fifoRdEntry <= "11";
                        o_RequestValid <= '1';
                    else -- Nothing available, go back to idle
                        rd_fsm <= idle;
                        o_RequestValid <= '0';
                    end if;
                    
                when waitRequest =>
                    if selectedPacketValid = '1' then
                        if (selectedOutputMux = OUTPUTMUX) then
                            rd_fsm <= sendData;
                        else
                            -- requested input port started to send something, but not to this output mux.
                            -- Go back to idle so we can try a different input port.
                            rd_fsm <= idle;
                        end if;
                    end if;
                
                when sendData =>
                    o_RequestValid <= '0';
                    if selectedPacketValid = '0' then
                        rd_fsm <= idle;
                    end if;
                
                when others =>
                    rd_fsm <= idle;
                    
            end case;
            
            rd_fsm_del <= rd_fsm;

            if rd_fsm = sendData and rd_fsm_del = waitRequest then
                fifoRd <= '1';
            else
                fifoRd <= '0';
            end if;
            
            selectedPacketValidDel <= selectedPacketValid;
            if ((selectedOutputMux = OUTPUTMUX) and (selectedPortPossible = '1')) then
                if DROPADDRWORD = '1' then
                    valid_int <= selectedPacketValid and selectedPacketValidDel;
                else
                    valid_int <= selectedPacketValid;
                end if;
            else
                valid_int <= '0';
            end if;
            o_data <= selectedPacketData;
            
            validDel <= valid_int;
            
            if rd_fsm = sendData and rd_fsm_del /= sendData and selectedPortPossible = '0' then
                oinputPortInvalid <= '1';
            else
                oinputPortInvalid <= '0';
            end if;
            
        end if;
    end process;
    o_valid <= valid_int;
    o_sop <= '1' when valid_int = '1' and validDel = '0' else '0';
    
    o_requestPort <= requestPort; -- The input port we are requesting data from.
    
    selectedPacketValid <= i_packetValid(to_integer(unsigned(requestPort)));
    selectedOutputMux <= i_packetOutputMux(to_integer(unsigned(requestPort)));
    selectedPortPossible <= PORTSUSED(to_integer(unsigned(requestPort)));
    
    maskGen: for i in 0 to 31 generate
        maskedPacketData(i) <= i_packetData(i) when PORTSUSED(i) = '1' else (others => '0');
    end generate;
    
    selectedPacketData <= maskedPacketData(to_integer(unsigned(requestPort)));
    
    process(i_IC_clk)
    begin
        if rising_edge(i_IC_clk) then
            if i_clrErrorCounts = '1' then
                anyPortInvalid <= '0';
                portInvalidCount <= "000";
                anyfifoFull <= '0';
                fifoFullCount <= "000";
            else
                if oinputPortInvalid = '1' then
                    anyPortInvalid <= '1';
                    portInvalidCount <= std_logic_vector(unsigned(portInvalidCount) + 1);
                end if;
                if ostatFifoFull = '1' then
                    anyfifoFull <= '1';
                    fifoFullCount <= std_logic_vector(unsigned(fifoFullCount) + 1);
                end if;
            end if;
        end if;
    end process;
    
    o_errCounts(3 downto 0) <= anyfifoFull & fifoFullCount;
    o_errCounts(7 downto 4) <= anyPortInvalid & portInvalidCount;
    
    
end Behavioral;

