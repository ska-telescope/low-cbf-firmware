LIBRARY IEEE, technology_lib;
USE IEEE.std_logic_1164.ALL;
USE technology_lib.technology_pkg.ALL;


PACKAGE tech_mac_40g_component_pkg IS

COMPONENT mac_40g_quad_122
  PORT (
    gt_rxp_in_0 : IN STD_LOGIC;
    gt_rxp_in_1 : IN STD_LOGIC;
    gt_rxp_in_2 : IN STD_LOGIC;
    gt_rxp_in_3 : IN STD_LOGIC;
    gt_rxn_in_0 : IN STD_LOGIC;
    gt_rxn_in_1 : IN STD_LOGIC;
    gt_rxn_in_2 : IN STD_LOGIC;
    gt_rxn_in_3 : IN STD_LOGIC;
    gt_txp_out_0 : OUT STD_LOGIC;
    gt_txp_out_1 : OUT STD_LOGIC;
    gt_txp_out_2 : OUT STD_LOGIC;
    gt_txp_out_3 : OUT STD_LOGIC;
    gt_txn_out_0 : OUT STD_LOGIC;
    gt_txn_out_1 : OUT STD_LOGIC;
    gt_txn_out_2 : OUT STD_LOGIC;
    gt_txn_out_3 : OUT STD_LOGIC;
    txoutclksel_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    rxoutclksel_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_dmonitorout_0 : OUT STD_LOGIC_VECTOR(67 DOWNTO 0);
    gt_eyescandataerror_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_eyescanreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_eyescantrigger_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_pcsrsvdin_0 : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
    gt_rxbufreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxbufstatus_0 : OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_rxcdrhold_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxcommadeten_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxdfeagchold_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxdfelpmreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxlatclk_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxlpmen_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpcsreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpmareset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpolarity_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbscntreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbserr_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbssel_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_rxrate_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_rxslide_in_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxstartofseq_0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    gt_txbufstatus_0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    gt_txdiffctrl_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gt_txinhibit_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txlatclk_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txmaincursor_0 : IN STD_LOGIC_VECTOR(27 DOWNTO 0);
    gt_txpcsreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpmareset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpolarity_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpostcursor_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gt_txprbsforceerr_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txprbssel_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_txprecursor_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gtwiz_reset_tx_datapath_0 : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    gtwiz_reset_rx_datapath_0 : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    rxrecclkout_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_common_drpclk : IN STD_LOGIC;
    gt_common_drpdo : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_common_drprdy : OUT STD_LOGIC;
    gt_common_drpen : IN STD_LOGIC;
    gt_common_drpwe : IN STD_LOGIC;
    gt_common_drpaddr : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_common_drpdi : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpclk_0 : IN STD_LOGIC;
    gt_ch_drpclk_1 : IN STD_LOGIC;
    gt_ch_drpclk_2 : IN STD_LOGIC;
    gt_ch_drpclk_3 : IN STD_LOGIC;
    gt_ch_drpdo_0 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_1 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_2 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_3 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drprdy_0 : OUT STD_LOGIC;
    gt_ch_drprdy_1 : OUT STD_LOGIC;
    gt_ch_drprdy_2 : OUT STD_LOGIC;
    gt_ch_drprdy_3 : OUT STD_LOGIC;
    gt_ch_drpen_0 : IN STD_LOGIC;
    gt_ch_drpen_1 : IN STD_LOGIC;
    gt_ch_drpen_2 : IN STD_LOGIC;
    gt_ch_drpen_3 : IN STD_LOGIC;
    gt_ch_drpwe_0 : IN STD_LOGIC;
    gt_ch_drpwe_1 : IN STD_LOGIC;
    gt_ch_drpwe_2 : IN STD_LOGIC;
    gt_ch_drpwe_3 : IN STD_LOGIC;
    gt_ch_drpaddr_0 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_1 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_2 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_3 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpdi_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_1 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_2 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_3 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    sys_reset : IN STD_LOGIC;
    dclk : IN STD_LOGIC;
    tx_clk_out_0 : OUT STD_LOGIC;
    rx_clk_out_0 : OUT STD_LOGIC;
    gt_refclk_p : IN STD_LOGIC;
    gt_refclk_n : IN STD_LOGIC;
    gt_refclk_out : OUT STD_LOGIC;
    gtpowergood_out_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    rx_reset_0 : IN STD_LOGIC;
    user_rx_reset_0 : OUT STD_LOGIC;
    rx_axis_tvalid_0 : OUT STD_LOGIC;
    rx_axis_tdata_0 : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
    rx_axis_tuser_0 : OUT STD_LOGIC_VECTOR(69 DOWNTO 0);
    ctl_rx_test_pattern_0 : IN STD_LOGIC;
    ctl_rx_enable_0 : IN STD_LOGIC;
    ctl_rx_delete_fcs_0 : IN STD_LOGIC;
    ctl_rx_ignore_fcs_0 : IN STD_LOGIC;
    ctl_rx_max_packet_len_0 : IN STD_LOGIC_VECTOR(14 DOWNTO 0);
    ctl_rx_min_packet_len_0 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    ctl_rx_custom_preamble_enable_0 : IN STD_LOGIC;
    ctl_rx_check_sfd_0 : IN STD_LOGIC;
    ctl_rx_check_preamble_0 : IN STD_LOGIC;
    ctl_rx_process_lfi_0 : IN STD_LOGIC;
    ctl_rx_force_resync_0 : IN STD_LOGIC;
    stat_rx_block_lock_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_framing_err_valid_0_0 : OUT STD_LOGIC;
    stat_rx_framing_err_0_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_1_0 : OUT STD_LOGIC;
    stat_rx_framing_err_1_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_2_0 : OUT STD_LOGIC;
    stat_rx_framing_err_2_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_3_0 : OUT STD_LOGIC;
    stat_rx_framing_err_3_0 : OUT STD_LOGIC;
    stat_rx_vl_demuxed_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_vl_number_0_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_1_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_2_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_3_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_synced_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_synced_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_len_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_repeat_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_misaligned_0 : OUT STD_LOGIC;
    stat_rx_aligned_err_0 : OUT STD_LOGIC;
    stat_rx_bip_err_0_0 : OUT STD_LOGIC;
    stat_rx_bip_err_1_0 : OUT STD_LOGIC;
    stat_rx_bip_err_2_0 : OUT STD_LOGIC;
    stat_rx_bip_err_3_0 : OUT STD_LOGIC;
    stat_rx_aligned_0 : OUT STD_LOGIC;
    stat_rx_hi_ber_0 : OUT STD_LOGIC;
    stat_rx_status_0 : OUT STD_LOGIC;
    stat_rx_bad_code_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_total_packets_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_total_good_packets_0 : OUT STD_LOGIC;
    stat_rx_total_bytes_0 : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    stat_rx_total_good_bytes_0 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_rx_packet_small_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_jabber_0 : OUT STD_LOGIC;
    stat_rx_packet_large_0 : OUT STD_LOGIC;
    stat_rx_oversize_0 : OUT STD_LOGIC;
    stat_rx_undersize_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_toolong_0 : OUT STD_LOGIC;
    stat_rx_fragment_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_64_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_65_127_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_128_255_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_256_511_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_512_1023_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1024_1518_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1519_1522_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1523_1548_bytes_0 : OUT STD_LOGIC;
    stat_rx_bad_fcs_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_bad_fcs_0 : OUT STD_LOGIC;
    stat_rx_stomped_fcs_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_1549_2047_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_2048_4095_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_4096_8191_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_8192_9215_bytes_0 : OUT STD_LOGIC;
    stat_rx_bad_preamble_0 : OUT STD_LOGIC;
    stat_rx_bad_sfd_0 : OUT STD_LOGIC;
    stat_rx_got_signal_os_0 : OUT STD_LOGIC;
    stat_rx_test_pattern_mismatch_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_truncated_0 : OUT STD_LOGIC;
    stat_rx_local_fault_0 : OUT STD_LOGIC;
    stat_rx_remote_fault_0 : OUT STD_LOGIC;
    stat_rx_internal_local_fault_0 : OUT STD_LOGIC;
    stat_rx_received_local_fault_0 : OUT STD_LOGIC;
    tx_reset_0 : IN STD_LOGIC;
    user_tx_reset_0 : OUT STD_LOGIC;
    tx_unfout_0 : OUT STD_LOGIC;
    tx_axis_tready_0 : OUT STD_LOGIC;
    tx_axis_tvalid_0 : IN STD_LOGIC;
    tx_axis_tdata_0 : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
    tx_axis_tuser_0 : IN STD_LOGIC_VECTOR(69 DOWNTO 0);
    stat_tx_total_packets_0 : OUT STD_LOGIC;
    stat_tx_total_bytes_0 : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
    stat_tx_total_good_packets_0 : OUT STD_LOGIC;
    stat_tx_total_good_bytes_0 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_tx_packet_64_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_65_127_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_128_255_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_256_511_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_512_1023_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1024_1518_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1519_1522_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1523_1548_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_small_0 : OUT STD_LOGIC;
    stat_tx_packet_large_0 : OUT STD_LOGIC;
    stat_tx_packet_1549_2047_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_2048_4095_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_4096_8191_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_8192_9215_bytes_0 : OUT STD_LOGIC;
    stat_tx_bad_fcs_0 : OUT STD_LOGIC;
    stat_tx_frame_error_0 : OUT STD_LOGIC;
    stat_tx_local_fault_0 : OUT STD_LOGIC;
    ctl_tx_test_pattern_0 : IN STD_LOGIC;
    ctl_tx_enable_0 : IN STD_LOGIC;
    ctl_tx_fcs_ins_enable_0 : IN STD_LOGIC;
    ctl_tx_ipg_value_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    ctl_tx_send_lfi_0 : IN STD_LOGIC;
    ctl_tx_send_rfi_0 : IN STD_LOGIC;
    ctl_tx_send_idle_0 : IN STD_LOGIC;
    ctl_tx_custom_preamble_enable_0 : IN STD_LOGIC;
    ctl_tx_ignore_fcs_0 : IN STD_LOGIC;
    gt_loopback_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    rx_core_clk_0 : IN STD_LOGIC
  );
END COMPONENT;

COMPONENT mac_40g_quad_124
  PORT (
    gt_rxp_in_0 : IN STD_LOGIC;
    gt_rxp_in_1 : IN STD_LOGIC;
    gt_rxp_in_2 : IN STD_LOGIC;
    gt_rxp_in_3 : IN STD_LOGIC;
    gt_rxn_in_0 : IN STD_LOGIC;
    gt_rxn_in_1 : IN STD_LOGIC;
    gt_rxn_in_2 : IN STD_LOGIC;
    gt_rxn_in_3 : IN STD_LOGIC;
    gt_txp_out_0 : OUT STD_LOGIC;
    gt_txp_out_1 : OUT STD_LOGIC;
    gt_txp_out_2 : OUT STD_LOGIC;
    gt_txp_out_3 : OUT STD_LOGIC;
    gt_txn_out_0 : OUT STD_LOGIC;
    gt_txn_out_1 : OUT STD_LOGIC;
    gt_txn_out_2 : OUT STD_LOGIC;
    gt_txn_out_3 : OUT STD_LOGIC;
    txoutclksel_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    rxoutclksel_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_dmonitorout_0 : OUT STD_LOGIC_VECTOR(67 DOWNTO 0);
    gt_eyescandataerror_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_eyescanreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_eyescantrigger_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_pcsrsvdin_0 : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
    gt_rxbufreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxbufstatus_0 : OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_rxcdrhold_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxcommadeten_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxdfeagchold_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxdfelpmreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxlatclk_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxlpmen_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpcsreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpmareset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpolarity_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbscntreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbserr_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbssel_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_rxrate_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_rxslide_in_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxstartofseq_0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    gt_txbufstatus_0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    gt_txdiffctrl_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gt_txinhibit_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txlatclk_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txmaincursor_0 : IN STD_LOGIC_VECTOR(27 DOWNTO 0);
    gt_txpcsreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpmareset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpolarity_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpostcursor_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gt_txprbsforceerr_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txprbssel_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_txprecursor_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gtwiz_reset_tx_datapath_0 : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    gtwiz_reset_rx_datapath_0 : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    rxrecclkout_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_common_drpclk : IN STD_LOGIC;
    gt_common_drpdo : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_common_drprdy : OUT STD_LOGIC;
    gt_common_drpen : IN STD_LOGIC;
    gt_common_drpwe : IN STD_LOGIC;
    gt_common_drpaddr : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_common_drpdi : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpclk_0 : IN STD_LOGIC;
    gt_ch_drpclk_1 : IN STD_LOGIC;
    gt_ch_drpclk_2 : IN STD_LOGIC;
    gt_ch_drpclk_3 : IN STD_LOGIC;
    gt_ch_drpdo_0 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_1 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_2 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_3 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drprdy_0 : OUT STD_LOGIC;
    gt_ch_drprdy_1 : OUT STD_LOGIC;
    gt_ch_drprdy_2 : OUT STD_LOGIC;
    gt_ch_drprdy_3 : OUT STD_LOGIC;
    gt_ch_drpen_0 : IN STD_LOGIC;
    gt_ch_drpen_1 : IN STD_LOGIC;
    gt_ch_drpen_2 : IN STD_LOGIC;
    gt_ch_drpen_3 : IN STD_LOGIC;
    gt_ch_drpwe_0 : IN STD_LOGIC;
    gt_ch_drpwe_1 : IN STD_LOGIC;
    gt_ch_drpwe_2 : IN STD_LOGIC;
    gt_ch_drpwe_3 : IN STD_LOGIC;
    gt_ch_drpaddr_0 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_1 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_2 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_3 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpdi_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_1 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_2 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_3 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    sys_reset : IN STD_LOGIC;
    dclk : IN STD_LOGIC;
    tx_clk_out_0 : OUT STD_LOGIC;
    rx_clk_out_0 : OUT STD_LOGIC;
    gt_refclk_p : IN STD_LOGIC;
    gt_refclk_n : IN STD_LOGIC;
    gt_refclk_out : OUT STD_LOGIC;
    gtpowergood_out_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    rx_reset_0 : IN STD_LOGIC;
    user_rx_reset_0 : OUT STD_LOGIC;
    rx_axis_tvalid_0 : OUT STD_LOGIC;
    rx_axis_tdata_0 : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
    rx_axis_tuser_0 : OUT STD_LOGIC_VECTOR(69 DOWNTO 0);
    ctl_rx_test_pattern_0 : IN STD_LOGIC;
    ctl_rx_enable_0 : IN STD_LOGIC;
    ctl_rx_delete_fcs_0 : IN STD_LOGIC;
    ctl_rx_ignore_fcs_0 : IN STD_LOGIC;
    ctl_rx_max_packet_len_0 : IN STD_LOGIC_VECTOR(14 DOWNTO 0);
    ctl_rx_min_packet_len_0 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    ctl_rx_custom_preamble_enable_0 : IN STD_LOGIC;
    ctl_rx_check_sfd_0 : IN STD_LOGIC;
    ctl_rx_check_preamble_0 : IN STD_LOGIC;
    ctl_rx_process_lfi_0 : IN STD_LOGIC;
    ctl_rx_force_resync_0 : IN STD_LOGIC;
    stat_rx_block_lock_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_framing_err_valid_0_0 : OUT STD_LOGIC;
    stat_rx_framing_err_0_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_1_0 : OUT STD_LOGIC;
    stat_rx_framing_err_1_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_2_0 : OUT STD_LOGIC;
    stat_rx_framing_err_2_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_3_0 : OUT STD_LOGIC;
    stat_rx_framing_err_3_0 : OUT STD_LOGIC;
    stat_rx_vl_demuxed_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_vl_number_0_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_1_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_2_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_3_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_synced_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_synced_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_len_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_repeat_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_misaligned_0 : OUT STD_LOGIC;
    stat_rx_aligned_err_0 : OUT STD_LOGIC;
    stat_rx_bip_err_0_0 : OUT STD_LOGIC;
    stat_rx_bip_err_1_0 : OUT STD_LOGIC;
    stat_rx_bip_err_2_0 : OUT STD_LOGIC;
    stat_rx_bip_err_3_0 : OUT STD_LOGIC;
    stat_rx_aligned_0 : OUT STD_LOGIC;
    stat_rx_hi_ber_0 : OUT STD_LOGIC;
    stat_rx_status_0 : OUT STD_LOGIC;
    stat_rx_bad_code_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_total_packets_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_total_good_packets_0 : OUT STD_LOGIC;
    stat_rx_total_bytes_0 : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    stat_rx_total_good_bytes_0 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_rx_packet_small_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_jabber_0 : OUT STD_LOGIC;
    stat_rx_packet_large_0 : OUT STD_LOGIC;
    stat_rx_oversize_0 : OUT STD_LOGIC;
    stat_rx_undersize_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_toolong_0 : OUT STD_LOGIC;
    stat_rx_fragment_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_64_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_65_127_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_128_255_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_256_511_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_512_1023_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1024_1518_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1519_1522_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1523_1548_bytes_0 : OUT STD_LOGIC;
    stat_rx_bad_fcs_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_bad_fcs_0 : OUT STD_LOGIC;
    stat_rx_stomped_fcs_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_1549_2047_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_2048_4095_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_4096_8191_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_8192_9215_bytes_0 : OUT STD_LOGIC;
    stat_rx_bad_preamble_0 : OUT STD_LOGIC;
    stat_rx_bad_sfd_0 : OUT STD_LOGIC;
    stat_rx_got_signal_os_0 : OUT STD_LOGIC;
    stat_rx_test_pattern_mismatch_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_truncated_0 : OUT STD_LOGIC;
    stat_rx_local_fault_0 : OUT STD_LOGIC;
    stat_rx_remote_fault_0 : OUT STD_LOGIC;
    stat_rx_internal_local_fault_0 : OUT STD_LOGIC;
    stat_rx_received_local_fault_0 : OUT STD_LOGIC;
    tx_reset_0 : IN STD_LOGIC;
    user_tx_reset_0 : OUT STD_LOGIC;
    tx_unfout_0 : OUT STD_LOGIC;
    tx_axis_tready_0 : OUT STD_LOGIC;
    tx_axis_tvalid_0 : IN STD_LOGIC;
    tx_axis_tdata_0 : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
    tx_axis_tuser_0 : IN STD_LOGIC_VECTOR(69 DOWNTO 0);
    stat_tx_total_packets_0 : OUT STD_LOGIC;
    stat_tx_total_bytes_0 : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
    stat_tx_total_good_packets_0 : OUT STD_LOGIC;
    stat_tx_total_good_bytes_0 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_tx_packet_64_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_65_127_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_128_255_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_256_511_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_512_1023_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1024_1518_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1519_1522_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1523_1548_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_small_0 : OUT STD_LOGIC;
    stat_tx_packet_large_0 : OUT STD_LOGIC;
    stat_tx_packet_1549_2047_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_2048_4095_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_4096_8191_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_8192_9215_bytes_0 : OUT STD_LOGIC;
    stat_tx_bad_fcs_0 : OUT STD_LOGIC;
    stat_tx_frame_error_0 : OUT STD_LOGIC;
    stat_tx_local_fault_0 : OUT STD_LOGIC;
    ctl_tx_test_pattern_0 : IN STD_LOGIC;
    ctl_tx_enable_0 : IN STD_LOGIC;
    ctl_tx_fcs_ins_enable_0 : IN STD_LOGIC;
    ctl_tx_ipg_value_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    ctl_tx_send_lfi_0 : IN STD_LOGIC;
    ctl_tx_send_rfi_0 : IN STD_LOGIC;
    ctl_tx_send_idle_0 : IN STD_LOGIC;
    ctl_tx_custom_preamble_enable_0 : IN STD_LOGIC;
    ctl_tx_ignore_fcs_0 : IN STD_LOGIC;
    gt_loopback_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    rx_core_clk_0 : IN STD_LOGIC
  );
END COMPONENT;

COMPONENT mac_40g_quad_125
  PORT (
    gt_rxp_in_0 : IN STD_LOGIC;
    gt_rxp_in_1 : IN STD_LOGIC;
    gt_rxp_in_2 : IN STD_LOGIC;
    gt_rxp_in_3 : IN STD_LOGIC;
    gt_rxn_in_0 : IN STD_LOGIC;
    gt_rxn_in_1 : IN STD_LOGIC;
    gt_rxn_in_2 : IN STD_LOGIC;
    gt_rxn_in_3 : IN STD_LOGIC;
    gt_txp_out_0 : OUT STD_LOGIC;
    gt_txp_out_1 : OUT STD_LOGIC;
    gt_txp_out_2 : OUT STD_LOGIC;
    gt_txp_out_3 : OUT STD_LOGIC;
    gt_txn_out_0 : OUT STD_LOGIC;
    gt_txn_out_1 : OUT STD_LOGIC;
    gt_txn_out_2 : OUT STD_LOGIC;
    gt_txn_out_3 : OUT STD_LOGIC;
    txoutclksel_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    rxoutclksel_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_dmonitorout_0 : OUT STD_LOGIC_VECTOR(67 DOWNTO 0);
    gt_eyescandataerror_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_eyescanreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_eyescantrigger_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_pcsrsvdin_0 : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
    gt_rxbufreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxbufstatus_0 : OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_rxcdrhold_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxcommadeten_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxdfeagchold_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxdfelpmreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxlatclk_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxlpmen_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpcsreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpmareset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpolarity_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbscntreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbserr_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbssel_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_rxrate_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_rxslide_in_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxstartofseq_0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    gt_txbufstatus_0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    gt_txdiffctrl_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gt_txinhibit_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txlatclk_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txmaincursor_0 : IN STD_LOGIC_VECTOR(27 DOWNTO 0);
    gt_txpcsreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpmareset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpolarity_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpostcursor_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gt_txprbsforceerr_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txprbssel_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_txprecursor_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gtwiz_reset_tx_datapath_0 : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    gtwiz_reset_rx_datapath_0 : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    rxrecclkout_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_common_drpclk : IN STD_LOGIC;
    gt_common_drpdo : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_common_drprdy : OUT STD_LOGIC;
    gt_common_drpen : IN STD_LOGIC;
    gt_common_drpwe : IN STD_LOGIC;
    gt_common_drpaddr : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_common_drpdi : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpclk_0 : IN STD_LOGIC;
    gt_ch_drpclk_1 : IN STD_LOGIC;
    gt_ch_drpclk_2 : IN STD_LOGIC;
    gt_ch_drpclk_3 : IN STD_LOGIC;
    gt_ch_drpdo_0 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_1 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_2 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_3 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drprdy_0 : OUT STD_LOGIC;
    gt_ch_drprdy_1 : OUT STD_LOGIC;
    gt_ch_drprdy_2 : OUT STD_LOGIC;
    gt_ch_drprdy_3 : OUT STD_LOGIC;
    gt_ch_drpen_0 : IN STD_LOGIC;
    gt_ch_drpen_1 : IN STD_LOGIC;
    gt_ch_drpen_2 : IN STD_LOGIC;
    gt_ch_drpen_3 : IN STD_LOGIC;
    gt_ch_drpwe_0 : IN STD_LOGIC;
    gt_ch_drpwe_1 : IN STD_LOGIC;
    gt_ch_drpwe_2 : IN STD_LOGIC;
    gt_ch_drpwe_3 : IN STD_LOGIC;
    gt_ch_drpaddr_0 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_1 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_2 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_3 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpdi_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_1 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_2 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_3 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    sys_reset : IN STD_LOGIC;
    dclk : IN STD_LOGIC;
    tx_clk_out_0 : OUT STD_LOGIC;
    rx_clk_out_0 : OUT STD_LOGIC;
    gt_refclk_p : IN STD_LOGIC;
    gt_refclk_n : IN STD_LOGIC;
    gt_refclk_out : OUT STD_LOGIC;
    gtpowergood_out_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    rx_reset_0 : IN STD_LOGIC;
    user_rx_reset_0 : OUT STD_LOGIC;
    rx_axis_tvalid_0 : OUT STD_LOGIC;
    rx_axis_tdata_0 : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
    rx_axis_tuser_0 : OUT STD_LOGIC_VECTOR(69 DOWNTO 0);
    ctl_rx_test_pattern_0 : IN STD_LOGIC;
    ctl_rx_enable_0 : IN STD_LOGIC;
    ctl_rx_delete_fcs_0 : IN STD_LOGIC;
    ctl_rx_ignore_fcs_0 : IN STD_LOGIC;
    ctl_rx_max_packet_len_0 : IN STD_LOGIC_VECTOR(14 DOWNTO 0);
    ctl_rx_min_packet_len_0 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    ctl_rx_custom_preamble_enable_0 : IN STD_LOGIC;
    ctl_rx_check_sfd_0 : IN STD_LOGIC;
    ctl_rx_check_preamble_0 : IN STD_LOGIC;
    ctl_rx_process_lfi_0 : IN STD_LOGIC;
    ctl_rx_force_resync_0 : IN STD_LOGIC;
    stat_rx_block_lock_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_framing_err_valid_0_0 : OUT STD_LOGIC;
    stat_rx_framing_err_0_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_1_0 : OUT STD_LOGIC;
    stat_rx_framing_err_1_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_2_0 : OUT STD_LOGIC;
    stat_rx_framing_err_2_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_3_0 : OUT STD_LOGIC;
    stat_rx_framing_err_3_0 : OUT STD_LOGIC;
    stat_rx_vl_demuxed_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_vl_number_0_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_1_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_2_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_3_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_synced_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_synced_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_len_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_repeat_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_misaligned_0 : OUT STD_LOGIC;
    stat_rx_aligned_err_0 : OUT STD_LOGIC;
    stat_rx_bip_err_0_0 : OUT STD_LOGIC;
    stat_rx_bip_err_1_0 : OUT STD_LOGIC;
    stat_rx_bip_err_2_0 : OUT STD_LOGIC;
    stat_rx_bip_err_3_0 : OUT STD_LOGIC;
    stat_rx_aligned_0 : OUT STD_LOGIC;
    stat_rx_hi_ber_0 : OUT STD_LOGIC;
    stat_rx_status_0 : OUT STD_LOGIC;
    stat_rx_bad_code_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_total_packets_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_total_good_packets_0 : OUT STD_LOGIC;
    stat_rx_total_bytes_0 : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    stat_rx_total_good_bytes_0 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_rx_packet_small_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_jabber_0 : OUT STD_LOGIC;
    stat_rx_packet_large_0 : OUT STD_LOGIC;
    stat_rx_oversize_0 : OUT STD_LOGIC;
    stat_rx_undersize_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_toolong_0 : OUT STD_LOGIC;
    stat_rx_fragment_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_64_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_65_127_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_128_255_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_256_511_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_512_1023_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1024_1518_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1519_1522_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1523_1548_bytes_0 : OUT STD_LOGIC;
    stat_rx_bad_fcs_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_bad_fcs_0 : OUT STD_LOGIC;
    stat_rx_stomped_fcs_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_1549_2047_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_2048_4095_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_4096_8191_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_8192_9215_bytes_0 : OUT STD_LOGIC;
    stat_rx_bad_preamble_0 : OUT STD_LOGIC;
    stat_rx_bad_sfd_0 : OUT STD_LOGIC;
    stat_rx_got_signal_os_0 : OUT STD_LOGIC;
    stat_rx_test_pattern_mismatch_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_truncated_0 : OUT STD_LOGIC;
    stat_rx_local_fault_0 : OUT STD_LOGIC;
    stat_rx_remote_fault_0 : OUT STD_LOGIC;
    stat_rx_internal_local_fault_0 : OUT STD_LOGIC;
    stat_rx_received_local_fault_0 : OUT STD_LOGIC;
    tx_reset_0 : IN STD_LOGIC;
    user_tx_reset_0 : OUT STD_LOGIC;
    tx_unfout_0 : OUT STD_LOGIC;
    tx_axis_tready_0 : OUT STD_LOGIC;
    tx_axis_tvalid_0 : IN STD_LOGIC;
    tx_axis_tdata_0 : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
    tx_axis_tuser_0 : IN STD_LOGIC_VECTOR(69 DOWNTO 0);
    stat_tx_total_packets_0 : OUT STD_LOGIC;
    stat_tx_total_bytes_0 : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
    stat_tx_total_good_packets_0 : OUT STD_LOGIC;
    stat_tx_total_good_bytes_0 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_tx_packet_64_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_65_127_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_128_255_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_256_511_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_512_1023_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1024_1518_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1519_1522_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1523_1548_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_small_0 : OUT STD_LOGIC;
    stat_tx_packet_large_0 : OUT STD_LOGIC;
    stat_tx_packet_1549_2047_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_2048_4095_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_4096_8191_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_8192_9215_bytes_0 : OUT STD_LOGIC;
    stat_tx_bad_fcs_0 : OUT STD_LOGIC;
    stat_tx_frame_error_0 : OUT STD_LOGIC;
    stat_tx_local_fault_0 : OUT STD_LOGIC;
    ctl_tx_test_pattern_0 : IN STD_LOGIC;
    ctl_tx_enable_0 : IN STD_LOGIC;
    ctl_tx_fcs_ins_enable_0 : IN STD_LOGIC;
    ctl_tx_ipg_value_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    ctl_tx_send_lfi_0 : IN STD_LOGIC;
    ctl_tx_send_rfi_0 : IN STD_LOGIC;
    ctl_tx_send_idle_0 : IN STD_LOGIC;
    ctl_tx_custom_preamble_enable_0 : IN STD_LOGIC;
    ctl_tx_ignore_fcs_0 : IN STD_LOGIC;
    gt_loopback_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    rx_core_clk_0 : IN STD_LOGIC
  );
END COMPONENT;

COMPONENT mac_40g_quad_126
  PORT (
    gt_rxp_in_0 : IN STD_LOGIC;
    gt_rxp_in_1 : IN STD_LOGIC;
    gt_rxp_in_2 : IN STD_LOGIC;
    gt_rxp_in_3 : IN STD_LOGIC;
    gt_rxn_in_0 : IN STD_LOGIC;
    gt_rxn_in_1 : IN STD_LOGIC;
    gt_rxn_in_2 : IN STD_LOGIC;
    gt_rxn_in_3 : IN STD_LOGIC;
    gt_txp_out_0 : OUT STD_LOGIC;
    gt_txp_out_1 : OUT STD_LOGIC;
    gt_txp_out_2 : OUT STD_LOGIC;
    gt_txp_out_3 : OUT STD_LOGIC;
    gt_txn_out_0 : OUT STD_LOGIC;
    gt_txn_out_1 : OUT STD_LOGIC;
    gt_txn_out_2 : OUT STD_LOGIC;
    gt_txn_out_3 : OUT STD_LOGIC;
    txoutclksel_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    rxoutclksel_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_dmonitorout_0 : OUT STD_LOGIC_VECTOR(67 DOWNTO 0);
    gt_eyescandataerror_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_eyescanreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_eyescantrigger_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_pcsrsvdin_0 : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
    gt_rxbufreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxbufstatus_0 : OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_rxcdrhold_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxcommadeten_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxdfeagchold_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxdfelpmreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxlatclk_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxlpmen_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpcsreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpmareset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpolarity_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbscntreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbserr_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbssel_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_rxrate_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_rxslide_in_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxstartofseq_0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    gt_txbufstatus_0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    gt_txdiffctrl_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gt_txinhibit_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txlatclk_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txmaincursor_0 : IN STD_LOGIC_VECTOR(27 DOWNTO 0);
    gt_txpcsreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpmareset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpolarity_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpostcursor_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gt_txprbsforceerr_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txprbssel_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_txprecursor_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gtwiz_reset_tx_datapath_0 : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    gtwiz_reset_rx_datapath_0 : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    rxrecclkout_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_common_drpclk : IN STD_LOGIC;
    gt_common_drpdo : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_common_drprdy : OUT STD_LOGIC;
    gt_common_drpen : IN STD_LOGIC;
    gt_common_drpwe : IN STD_LOGIC;
    gt_common_drpaddr : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_common_drpdi : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpclk_0 : IN STD_LOGIC;
    gt_ch_drpclk_1 : IN STD_LOGIC;
    gt_ch_drpclk_2 : IN STD_LOGIC;
    gt_ch_drpclk_3 : IN STD_LOGIC;
    gt_ch_drpdo_0 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_1 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_2 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_3 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drprdy_0 : OUT STD_LOGIC;
    gt_ch_drprdy_1 : OUT STD_LOGIC;
    gt_ch_drprdy_2 : OUT STD_LOGIC;
    gt_ch_drprdy_3 : OUT STD_LOGIC;
    gt_ch_drpen_0 : IN STD_LOGIC;
    gt_ch_drpen_1 : IN STD_LOGIC;
    gt_ch_drpen_2 : IN STD_LOGIC;
    gt_ch_drpen_3 : IN STD_LOGIC;
    gt_ch_drpwe_0 : IN STD_LOGIC;
    gt_ch_drpwe_1 : IN STD_LOGIC;
    gt_ch_drpwe_2 : IN STD_LOGIC;
    gt_ch_drpwe_3 : IN STD_LOGIC;
    gt_ch_drpaddr_0 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_1 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_2 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_3 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpdi_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_1 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_2 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_3 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    sys_reset : IN STD_LOGIC;
    dclk : IN STD_LOGIC;
    tx_clk_out_0 : OUT STD_LOGIC;
    rx_clk_out_0 : OUT STD_LOGIC;
    gt_refclk_p : IN STD_LOGIC;
    gt_refclk_n : IN STD_LOGIC;
    gt_refclk_out : OUT STD_LOGIC;
    gtpowergood_out_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    rx_reset_0 : IN STD_LOGIC;
    user_rx_reset_0 : OUT STD_LOGIC;
    rx_axis_tvalid_0 : OUT STD_LOGIC;
    rx_axis_tdata_0 : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
    rx_axis_tuser_0 : OUT STD_LOGIC_VECTOR(69 DOWNTO 0);
    ctl_rx_test_pattern_0 : IN STD_LOGIC;
    ctl_rx_enable_0 : IN STD_LOGIC;
    ctl_rx_delete_fcs_0 : IN STD_LOGIC;
    ctl_rx_ignore_fcs_0 : IN STD_LOGIC;
    ctl_rx_max_packet_len_0 : IN STD_LOGIC_VECTOR(14 DOWNTO 0);
    ctl_rx_min_packet_len_0 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    ctl_rx_custom_preamble_enable_0 : IN STD_LOGIC;
    ctl_rx_check_sfd_0 : IN STD_LOGIC;
    ctl_rx_check_preamble_0 : IN STD_LOGIC;
    ctl_rx_process_lfi_0 : IN STD_LOGIC;
    ctl_rx_force_resync_0 : IN STD_LOGIC;
    stat_rx_block_lock_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_framing_err_valid_0_0 : OUT STD_LOGIC;
    stat_rx_framing_err_0_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_1_0 : OUT STD_LOGIC;
    stat_rx_framing_err_1_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_2_0 : OUT STD_LOGIC;
    stat_rx_framing_err_2_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_3_0 : OUT STD_LOGIC;
    stat_rx_framing_err_3_0 : OUT STD_LOGIC;
    stat_rx_vl_demuxed_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_vl_number_0_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_1_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_2_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_3_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_synced_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_synced_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_len_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_repeat_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_misaligned_0 : OUT STD_LOGIC;
    stat_rx_aligned_err_0 : OUT STD_LOGIC;
    stat_rx_bip_err_0_0 : OUT STD_LOGIC;
    stat_rx_bip_err_1_0 : OUT STD_LOGIC;
    stat_rx_bip_err_2_0 : OUT STD_LOGIC;
    stat_rx_bip_err_3_0 : OUT STD_LOGIC;
    stat_rx_aligned_0 : OUT STD_LOGIC;
    stat_rx_hi_ber_0 : OUT STD_LOGIC;
    stat_rx_status_0 : OUT STD_LOGIC;
    stat_rx_bad_code_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_total_packets_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_total_good_packets_0 : OUT STD_LOGIC;
    stat_rx_total_bytes_0 : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    stat_rx_total_good_bytes_0 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_rx_packet_small_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_jabber_0 : OUT STD_LOGIC;
    stat_rx_packet_large_0 : OUT STD_LOGIC;
    stat_rx_oversize_0 : OUT STD_LOGIC;
    stat_rx_undersize_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_toolong_0 : OUT STD_LOGIC;
    stat_rx_fragment_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_64_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_65_127_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_128_255_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_256_511_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_512_1023_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1024_1518_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1519_1522_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1523_1548_bytes_0 : OUT STD_LOGIC;
    stat_rx_bad_fcs_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_bad_fcs_0 : OUT STD_LOGIC;
    stat_rx_stomped_fcs_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_1549_2047_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_2048_4095_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_4096_8191_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_8192_9215_bytes_0 : OUT STD_LOGIC;
    stat_rx_bad_preamble_0 : OUT STD_LOGIC;
    stat_rx_bad_sfd_0 : OUT STD_LOGIC;
    stat_rx_got_signal_os_0 : OUT STD_LOGIC;
    stat_rx_test_pattern_mismatch_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_truncated_0 : OUT STD_LOGIC;
    stat_rx_local_fault_0 : OUT STD_LOGIC;
    stat_rx_remote_fault_0 : OUT STD_LOGIC;
    stat_rx_internal_local_fault_0 : OUT STD_LOGIC;
    stat_rx_received_local_fault_0 : OUT STD_LOGIC;
    tx_reset_0 : IN STD_LOGIC;
    user_tx_reset_0 : OUT STD_LOGIC;
    tx_unfout_0 : OUT STD_LOGIC;
    tx_axis_tready_0 : OUT STD_LOGIC;
    tx_axis_tvalid_0 : IN STD_LOGIC;
    tx_axis_tdata_0 : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
    tx_axis_tuser_0 : IN STD_LOGIC_VECTOR(69 DOWNTO 0);
    stat_tx_total_packets_0 : OUT STD_LOGIC;
    stat_tx_total_bytes_0 : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
    stat_tx_total_good_packets_0 : OUT STD_LOGIC;
    stat_tx_total_good_bytes_0 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_tx_packet_64_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_65_127_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_128_255_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_256_511_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_512_1023_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1024_1518_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1519_1522_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1523_1548_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_small_0 : OUT STD_LOGIC;
    stat_tx_packet_large_0 : OUT STD_LOGIC;
    stat_tx_packet_1549_2047_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_2048_4095_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_4096_8191_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_8192_9215_bytes_0 : OUT STD_LOGIC;
    stat_tx_bad_fcs_0 : OUT STD_LOGIC;
    stat_tx_frame_error_0 : OUT STD_LOGIC;
    stat_tx_local_fault_0 : OUT STD_LOGIC;
    ctl_tx_test_pattern_0 : IN STD_LOGIC;
    ctl_tx_enable_0 : IN STD_LOGIC;
    ctl_tx_fcs_ins_enable_0 : IN STD_LOGIC;
    ctl_tx_ipg_value_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    ctl_tx_send_lfi_0 : IN STD_LOGIC;
    ctl_tx_send_rfi_0 : IN STD_LOGIC;
    ctl_tx_send_idle_0 : IN STD_LOGIC;
    ctl_tx_custom_preamble_enable_0 : IN STD_LOGIC;
    ctl_tx_ignore_fcs_0 : IN STD_LOGIC;
    gt_loopback_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    rx_core_clk_0 : IN STD_LOGIC
  );
END COMPONENT;

COMPONENT mac_40g_quad_128
  PORT (
    gt_rxp_in_0 : IN STD_LOGIC;
    gt_rxp_in_1 : IN STD_LOGIC;
    gt_rxp_in_2 : IN STD_LOGIC;
    gt_rxp_in_3 : IN STD_LOGIC;
    gt_rxn_in_0 : IN STD_LOGIC;
    gt_rxn_in_1 : IN STD_LOGIC;
    gt_rxn_in_2 : IN STD_LOGIC;
    gt_rxn_in_3 : IN STD_LOGIC;
    gt_txp_out_0 : OUT STD_LOGIC;
    gt_txp_out_1 : OUT STD_LOGIC;
    gt_txp_out_2 : OUT STD_LOGIC;
    gt_txp_out_3 : OUT STD_LOGIC;
    gt_txn_out_0 : OUT STD_LOGIC;
    gt_txn_out_1 : OUT STD_LOGIC;
    gt_txn_out_2 : OUT STD_LOGIC;
    gt_txn_out_3 : OUT STD_LOGIC;
    txoutclksel_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    rxoutclksel_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_dmonitorout_0 : OUT STD_LOGIC_VECTOR(67 DOWNTO 0);
    gt_eyescandataerror_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_eyescanreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_eyescantrigger_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_pcsrsvdin_0 : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
    gt_rxbufreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxbufstatus_0 : OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_rxcdrhold_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxcommadeten_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxdfeagchold_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxdfelpmreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxlatclk_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxlpmen_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpcsreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpmareset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpolarity_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbscntreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbserr_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbssel_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_rxrate_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_rxslide_in_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxstartofseq_0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    gt_txbufstatus_0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    gt_txdiffctrl_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gt_txinhibit_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txlatclk_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txmaincursor_0 : IN STD_LOGIC_VECTOR(27 DOWNTO 0);
    gt_txpcsreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpmareset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpolarity_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpostcursor_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gt_txprbsforceerr_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txprbssel_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_txprecursor_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gtwiz_reset_tx_datapath_0 : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    gtwiz_reset_rx_datapath_0 : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    rxrecclkout_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_common_drpclk : IN STD_LOGIC;
    gt_common_drpdo : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_common_drprdy : OUT STD_LOGIC;
    gt_common_drpen : IN STD_LOGIC;
    gt_common_drpwe : IN STD_LOGIC;
    gt_common_drpaddr : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_common_drpdi : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpclk_0 : IN STD_LOGIC;
    gt_ch_drpclk_1 : IN STD_LOGIC;
    gt_ch_drpclk_2 : IN STD_LOGIC;
    gt_ch_drpclk_3 : IN STD_LOGIC;
    gt_ch_drpdo_0 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_1 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_2 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_3 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drprdy_0 : OUT STD_LOGIC;
    gt_ch_drprdy_1 : OUT STD_LOGIC;
    gt_ch_drprdy_2 : OUT STD_LOGIC;
    gt_ch_drprdy_3 : OUT STD_LOGIC;
    gt_ch_drpen_0 : IN STD_LOGIC;
    gt_ch_drpen_1 : IN STD_LOGIC;
    gt_ch_drpen_2 : IN STD_LOGIC;
    gt_ch_drpen_3 : IN STD_LOGIC;
    gt_ch_drpwe_0 : IN STD_LOGIC;
    gt_ch_drpwe_1 : IN STD_LOGIC;
    gt_ch_drpwe_2 : IN STD_LOGIC;
    gt_ch_drpwe_3 : IN STD_LOGIC;
    gt_ch_drpaddr_0 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_1 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_2 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_3 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpdi_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_1 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_2 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_3 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    sys_reset : IN STD_LOGIC;
    dclk : IN STD_LOGIC;
    tx_clk_out_0 : OUT STD_LOGIC;
    rx_clk_out_0 : OUT STD_LOGIC;
    gt_refclk_p : IN STD_LOGIC;
    gt_refclk_n : IN STD_LOGIC;
    gt_refclk_out : OUT STD_LOGIC;
    gtpowergood_out_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    rx_reset_0 : IN STD_LOGIC;
    user_rx_reset_0 : OUT STD_LOGIC;
    rx_axis_tvalid_0 : OUT STD_LOGIC;
    rx_axis_tdata_0 : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
    rx_axis_tuser_0 : OUT STD_LOGIC_VECTOR(69 DOWNTO 0);
    ctl_rx_test_pattern_0 : IN STD_LOGIC;
    ctl_rx_enable_0 : IN STD_LOGIC;
    ctl_rx_delete_fcs_0 : IN STD_LOGIC;
    ctl_rx_ignore_fcs_0 : IN STD_LOGIC;
    ctl_rx_max_packet_len_0 : IN STD_LOGIC_VECTOR(14 DOWNTO 0);
    ctl_rx_min_packet_len_0 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    ctl_rx_custom_preamble_enable_0 : IN STD_LOGIC;
    ctl_rx_check_sfd_0 : IN STD_LOGIC;
    ctl_rx_check_preamble_0 : IN STD_LOGIC;
    ctl_rx_process_lfi_0 : IN STD_LOGIC;
    ctl_rx_force_resync_0 : IN STD_LOGIC;
    stat_rx_block_lock_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_framing_err_valid_0_0 : OUT STD_LOGIC;
    stat_rx_framing_err_0_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_1_0 : OUT STD_LOGIC;
    stat_rx_framing_err_1_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_2_0 : OUT STD_LOGIC;
    stat_rx_framing_err_2_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_3_0 : OUT STD_LOGIC;
    stat_rx_framing_err_3_0 : OUT STD_LOGIC;
    stat_rx_vl_demuxed_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_vl_number_0_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_1_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_2_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_3_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_synced_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_synced_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_len_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_repeat_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_misaligned_0 : OUT STD_LOGIC;
    stat_rx_aligned_err_0 : OUT STD_LOGIC;
    stat_rx_bip_err_0_0 : OUT STD_LOGIC;
    stat_rx_bip_err_1_0 : OUT STD_LOGIC;
    stat_rx_bip_err_2_0 : OUT STD_LOGIC;
    stat_rx_bip_err_3_0 : OUT STD_LOGIC;
    stat_rx_aligned_0 : OUT STD_LOGIC;
    stat_rx_hi_ber_0 : OUT STD_LOGIC;
    stat_rx_status_0 : OUT STD_LOGIC;
    stat_rx_bad_code_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_total_packets_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_total_good_packets_0 : OUT STD_LOGIC;
    stat_rx_total_bytes_0 : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    stat_rx_total_good_bytes_0 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_rx_packet_small_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_jabber_0 : OUT STD_LOGIC;
    stat_rx_packet_large_0 : OUT STD_LOGIC;
    stat_rx_oversize_0 : OUT STD_LOGIC;
    stat_rx_undersize_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_toolong_0 : OUT STD_LOGIC;
    stat_rx_fragment_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_64_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_65_127_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_128_255_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_256_511_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_512_1023_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1024_1518_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1519_1522_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1523_1548_bytes_0 : OUT STD_LOGIC;
    stat_rx_bad_fcs_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_bad_fcs_0 : OUT STD_LOGIC;
    stat_rx_stomped_fcs_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_1549_2047_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_2048_4095_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_4096_8191_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_8192_9215_bytes_0 : OUT STD_LOGIC;
    stat_rx_bad_preamble_0 : OUT STD_LOGIC;
    stat_rx_bad_sfd_0 : OUT STD_LOGIC;
    stat_rx_got_signal_os_0 : OUT STD_LOGIC;
    stat_rx_test_pattern_mismatch_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_truncated_0 : OUT STD_LOGIC;
    stat_rx_local_fault_0 : OUT STD_LOGIC;
    stat_rx_remote_fault_0 : OUT STD_LOGIC;
    stat_rx_internal_local_fault_0 : OUT STD_LOGIC;
    stat_rx_received_local_fault_0 : OUT STD_LOGIC;
    tx_reset_0 : IN STD_LOGIC;
    user_tx_reset_0 : OUT STD_LOGIC;
    tx_unfout_0 : OUT STD_LOGIC;
    tx_axis_tready_0 : OUT STD_LOGIC;
    tx_axis_tvalid_0 : IN STD_LOGIC;
    tx_axis_tdata_0 : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
    tx_axis_tuser_0 : IN STD_LOGIC_VECTOR(69 DOWNTO 0);
    stat_tx_total_packets_0 : OUT STD_LOGIC;
    stat_tx_total_bytes_0 : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
    stat_tx_total_good_packets_0 : OUT STD_LOGIC;
    stat_tx_total_good_bytes_0 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_tx_packet_64_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_65_127_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_128_255_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_256_511_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_512_1023_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1024_1518_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1519_1522_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1523_1548_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_small_0 : OUT STD_LOGIC;
    stat_tx_packet_large_0 : OUT STD_LOGIC;
    stat_tx_packet_1549_2047_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_2048_4095_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_4096_8191_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_8192_9215_bytes_0 : OUT STD_LOGIC;
    stat_tx_bad_fcs_0 : OUT STD_LOGIC;
    stat_tx_frame_error_0 : OUT STD_LOGIC;
    stat_tx_local_fault_0 : OUT STD_LOGIC;
    ctl_tx_test_pattern_0 : IN STD_LOGIC;
    ctl_tx_enable_0 : IN STD_LOGIC;
    ctl_tx_fcs_ins_enable_0 : IN STD_LOGIC;
    ctl_tx_ipg_value_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    ctl_tx_send_lfi_0 : IN STD_LOGIC;
    ctl_tx_send_rfi_0 : IN STD_LOGIC;
    ctl_tx_send_idle_0 : IN STD_LOGIC;
    ctl_tx_custom_preamble_enable_0 : IN STD_LOGIC;
    ctl_tx_ignore_fcs_0 : IN STD_LOGIC;
    gt_loopback_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    rx_core_clk_0 : IN STD_LOGIC
  );
END COMPONENT;

COMPONENT mac_40g_quad_130
  PORT (
    gt_rxp_in_0 : IN STD_LOGIC;
    gt_rxp_in_1 : IN STD_LOGIC;
    gt_rxp_in_2 : IN STD_LOGIC;
    gt_rxp_in_3 : IN STD_LOGIC;
    gt_rxn_in_0 : IN STD_LOGIC;
    gt_rxn_in_1 : IN STD_LOGIC;
    gt_rxn_in_2 : IN STD_LOGIC;
    gt_rxn_in_3 : IN STD_LOGIC;
    gt_txp_out_0 : OUT STD_LOGIC;
    gt_txp_out_1 : OUT STD_LOGIC;
    gt_txp_out_2 : OUT STD_LOGIC;
    gt_txp_out_3 : OUT STD_LOGIC;
    gt_txn_out_0 : OUT STD_LOGIC;
    gt_txn_out_1 : OUT STD_LOGIC;
    gt_txn_out_2 : OUT STD_LOGIC;
    gt_txn_out_3 : OUT STD_LOGIC;
    txoutclksel_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    rxoutclksel_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_dmonitorout_0 : OUT STD_LOGIC_VECTOR(67 DOWNTO 0);
    gt_eyescandataerror_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_eyescanreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_eyescantrigger_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_pcsrsvdin_0 : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
    gt_rxbufreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxbufstatus_0 : OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_rxcdrhold_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxcommadeten_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxdfeagchold_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxdfelpmreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxlatclk_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxlpmen_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpcsreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpmareset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpolarity_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbscntreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbserr_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbssel_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_rxrate_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_rxslide_in_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxstartofseq_0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    gt_txbufstatus_0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    gt_txdiffctrl_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gt_txinhibit_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txlatclk_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txmaincursor_0 : IN STD_LOGIC_VECTOR(27 DOWNTO 0);
    gt_txpcsreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpmareset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpolarity_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpostcursor_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gt_txprbsforceerr_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txprbssel_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_txprecursor_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gtwiz_reset_tx_datapath_0 : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    gtwiz_reset_rx_datapath_0 : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    rxrecclkout_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_common_drpclk : IN STD_LOGIC;
    gt_common_drpdo : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_common_drprdy : OUT STD_LOGIC;
    gt_common_drpen : IN STD_LOGIC;
    gt_common_drpwe : IN STD_LOGIC;
    gt_common_drpaddr : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_common_drpdi : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpclk_0 : IN STD_LOGIC;
    gt_ch_drpclk_1 : IN STD_LOGIC;
    gt_ch_drpclk_2 : IN STD_LOGIC;
    gt_ch_drpclk_3 : IN STD_LOGIC;
    gt_ch_drpdo_0 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_1 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_2 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_3 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drprdy_0 : OUT STD_LOGIC;
    gt_ch_drprdy_1 : OUT STD_LOGIC;
    gt_ch_drprdy_2 : OUT STD_LOGIC;
    gt_ch_drprdy_3 : OUT STD_LOGIC;
    gt_ch_drpen_0 : IN STD_LOGIC;
    gt_ch_drpen_1 : IN STD_LOGIC;
    gt_ch_drpen_2 : IN STD_LOGIC;
    gt_ch_drpen_3 : IN STD_LOGIC;
    gt_ch_drpwe_0 : IN STD_LOGIC;
    gt_ch_drpwe_1 : IN STD_LOGIC;
    gt_ch_drpwe_2 : IN STD_LOGIC;
    gt_ch_drpwe_3 : IN STD_LOGIC;
    gt_ch_drpaddr_0 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_1 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_2 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_3 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpdi_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_1 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_2 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_3 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    sys_reset : IN STD_LOGIC;
    dclk : IN STD_LOGIC;
    tx_clk_out_0 : OUT STD_LOGIC;
    rx_clk_out_0 : OUT STD_LOGIC;
    gt_refclk_p : IN STD_LOGIC;
    gt_refclk_n : IN STD_LOGIC;
    gt_refclk_out : OUT STD_LOGIC;
    gtpowergood_out_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    rx_reset_0 : IN STD_LOGIC;
    user_rx_reset_0 : OUT STD_LOGIC;
    rx_axis_tvalid_0 : OUT STD_LOGIC;
    rx_axis_tdata_0 : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
    rx_axis_tuser_0 : OUT STD_LOGIC_VECTOR(69 DOWNTO 0);
    ctl_rx_test_pattern_0 : IN STD_LOGIC;
    ctl_rx_enable_0 : IN STD_LOGIC;
    ctl_rx_delete_fcs_0 : IN STD_LOGIC;
    ctl_rx_ignore_fcs_0 : IN STD_LOGIC;
    ctl_rx_max_packet_len_0 : IN STD_LOGIC_VECTOR(14 DOWNTO 0);
    ctl_rx_min_packet_len_0 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    ctl_rx_custom_preamble_enable_0 : IN STD_LOGIC;
    ctl_rx_check_sfd_0 : IN STD_LOGIC;
    ctl_rx_check_preamble_0 : IN STD_LOGIC;
    ctl_rx_process_lfi_0 : IN STD_LOGIC;
    ctl_rx_force_resync_0 : IN STD_LOGIC;
    stat_rx_block_lock_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_framing_err_valid_0_0 : OUT STD_LOGIC;
    stat_rx_framing_err_0_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_1_0 : OUT STD_LOGIC;
    stat_rx_framing_err_1_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_2_0 : OUT STD_LOGIC;
    stat_rx_framing_err_2_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_3_0 : OUT STD_LOGIC;
    stat_rx_framing_err_3_0 : OUT STD_LOGIC;
    stat_rx_vl_demuxed_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_vl_number_0_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_1_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_2_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_3_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_synced_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_synced_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_len_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_repeat_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_misaligned_0 : OUT STD_LOGIC;
    stat_rx_aligned_err_0 : OUT STD_LOGIC;
    stat_rx_bip_err_0_0 : OUT STD_LOGIC;
    stat_rx_bip_err_1_0 : OUT STD_LOGIC;
    stat_rx_bip_err_2_0 : OUT STD_LOGIC;
    stat_rx_bip_err_3_0 : OUT STD_LOGIC;
    stat_rx_aligned_0 : OUT STD_LOGIC;
    stat_rx_hi_ber_0 : OUT STD_LOGIC;
    stat_rx_status_0 : OUT STD_LOGIC;
    stat_rx_bad_code_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_total_packets_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_total_good_packets_0 : OUT STD_LOGIC;
    stat_rx_total_bytes_0 : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    stat_rx_total_good_bytes_0 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_rx_packet_small_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_jabber_0 : OUT STD_LOGIC;
    stat_rx_packet_large_0 : OUT STD_LOGIC;
    stat_rx_oversize_0 : OUT STD_LOGIC;
    stat_rx_undersize_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_toolong_0 : OUT STD_LOGIC;
    stat_rx_fragment_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_64_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_65_127_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_128_255_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_256_511_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_512_1023_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1024_1518_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1519_1522_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1523_1548_bytes_0 : OUT STD_LOGIC;
    stat_rx_bad_fcs_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_bad_fcs_0 : OUT STD_LOGIC;
    stat_rx_stomped_fcs_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_1549_2047_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_2048_4095_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_4096_8191_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_8192_9215_bytes_0 : OUT STD_LOGIC;
    stat_rx_bad_preamble_0 : OUT STD_LOGIC;
    stat_rx_bad_sfd_0 : OUT STD_LOGIC;
    stat_rx_got_signal_os_0 : OUT STD_LOGIC;
    stat_rx_test_pattern_mismatch_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_truncated_0 : OUT STD_LOGIC;
    stat_rx_local_fault_0 : OUT STD_LOGIC;
    stat_rx_remote_fault_0 : OUT STD_LOGIC;
    stat_rx_internal_local_fault_0 : OUT STD_LOGIC;
    stat_rx_received_local_fault_0 : OUT STD_LOGIC;
    tx_reset_0 : IN STD_LOGIC;
    user_tx_reset_0 : OUT STD_LOGIC;
    tx_unfout_0 : OUT STD_LOGIC;
    tx_axis_tready_0 : OUT STD_LOGIC;
    tx_axis_tvalid_0 : IN STD_LOGIC;
    tx_axis_tdata_0 : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
    tx_axis_tuser_0 : IN STD_LOGIC_VECTOR(69 DOWNTO 0);
    stat_tx_total_packets_0 : OUT STD_LOGIC;
    stat_tx_total_bytes_0 : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
    stat_tx_total_good_packets_0 : OUT STD_LOGIC;
    stat_tx_total_good_bytes_0 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_tx_packet_64_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_65_127_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_128_255_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_256_511_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_512_1023_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1024_1518_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1519_1522_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1523_1548_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_small_0 : OUT STD_LOGIC;
    stat_tx_packet_large_0 : OUT STD_LOGIC;
    stat_tx_packet_1549_2047_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_2048_4095_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_4096_8191_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_8192_9215_bytes_0 : OUT STD_LOGIC;
    stat_tx_bad_fcs_0 : OUT STD_LOGIC;
    stat_tx_frame_error_0 : OUT STD_LOGIC;
    stat_tx_local_fault_0 : OUT STD_LOGIC;
    ctl_tx_test_pattern_0 : IN STD_LOGIC;
    ctl_tx_enable_0 : IN STD_LOGIC;
    ctl_tx_fcs_ins_enable_0 : IN STD_LOGIC;
    ctl_tx_ipg_value_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    ctl_tx_send_lfi_0 : IN STD_LOGIC;
    ctl_tx_send_rfi_0 : IN STD_LOGIC;
    ctl_tx_send_idle_0 : IN STD_LOGIC;
    ctl_tx_custom_preamble_enable_0 : IN STD_LOGIC;
    ctl_tx_ignore_fcs_0 : IN STD_LOGIC;
    gt_loopback_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    rx_core_clk_0 : IN STD_LOGIC
  );
END COMPONENT;

COMPONENT mac_40g_quad_131
  PORT (
    gt_rxp_in_0 : IN STD_LOGIC;
    gt_rxp_in_1 : IN STD_LOGIC;
    gt_rxp_in_2 : IN STD_LOGIC;
    gt_rxp_in_3 : IN STD_LOGIC;
    gt_rxn_in_0 : IN STD_LOGIC;
    gt_rxn_in_1 : IN STD_LOGIC;
    gt_rxn_in_2 : IN STD_LOGIC;
    gt_rxn_in_3 : IN STD_LOGIC;
    gt_txp_out_0 : OUT STD_LOGIC;
    gt_txp_out_1 : OUT STD_LOGIC;
    gt_txp_out_2 : OUT STD_LOGIC;
    gt_txp_out_3 : OUT STD_LOGIC;
    gt_txn_out_0 : OUT STD_LOGIC;
    gt_txn_out_1 : OUT STD_LOGIC;
    gt_txn_out_2 : OUT STD_LOGIC;
    gt_txn_out_3 : OUT STD_LOGIC;
    txoutclksel_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    rxoutclksel_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_dmonitorout_0 : OUT STD_LOGIC_VECTOR(67 DOWNTO 0);
    gt_eyescandataerror_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_eyescanreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_eyescantrigger_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_pcsrsvdin_0 : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
    gt_rxbufreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxbufstatus_0 : OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_rxcdrhold_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxcommadeten_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxdfeagchold_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxdfelpmreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxlatclk_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxlpmen_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpcsreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpmareset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpolarity_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbscntreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbserr_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbssel_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_rxrate_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_rxslide_in_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxstartofseq_0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    gt_txbufstatus_0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    gt_txdiffctrl_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gt_txinhibit_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txlatclk_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txmaincursor_0 : IN STD_LOGIC_VECTOR(27 DOWNTO 0);
    gt_txpcsreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpmareset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpolarity_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpostcursor_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gt_txprbsforceerr_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txprbssel_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_txprecursor_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gtwiz_reset_tx_datapath_0 : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    gtwiz_reset_rx_datapath_0 : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    rxrecclkout_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_common_drpclk : IN STD_LOGIC;
    gt_common_drpdo : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_common_drprdy : OUT STD_LOGIC;
    gt_common_drpen : IN STD_LOGIC;
    gt_common_drpwe : IN STD_LOGIC;
    gt_common_drpaddr : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_common_drpdi : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpclk_0 : IN STD_LOGIC;
    gt_ch_drpclk_1 : IN STD_LOGIC;
    gt_ch_drpclk_2 : IN STD_LOGIC;
    gt_ch_drpclk_3 : IN STD_LOGIC;
    gt_ch_drpdo_0 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_1 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_2 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_3 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drprdy_0 : OUT STD_LOGIC;
    gt_ch_drprdy_1 : OUT STD_LOGIC;
    gt_ch_drprdy_2 : OUT STD_LOGIC;
    gt_ch_drprdy_3 : OUT STD_LOGIC;
    gt_ch_drpen_0 : IN STD_LOGIC;
    gt_ch_drpen_1 : IN STD_LOGIC;
    gt_ch_drpen_2 : IN STD_LOGIC;
    gt_ch_drpen_3 : IN STD_LOGIC;
    gt_ch_drpwe_0 : IN STD_LOGIC;
    gt_ch_drpwe_1 : IN STD_LOGIC;
    gt_ch_drpwe_2 : IN STD_LOGIC;
    gt_ch_drpwe_3 : IN STD_LOGIC;
    gt_ch_drpaddr_0 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_1 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_2 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_3 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpdi_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_1 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_2 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_3 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    sys_reset : IN STD_LOGIC;
    dclk : IN STD_LOGIC;
    tx_clk_out_0 : OUT STD_LOGIC;
    rx_clk_out_0 : OUT STD_LOGIC;
    gt_refclk_p : IN STD_LOGIC;
    gt_refclk_n : IN STD_LOGIC;
    gt_refclk_out : OUT STD_LOGIC;
    gtpowergood_out_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    rx_reset_0 : IN STD_LOGIC;
    user_rx_reset_0 : OUT STD_LOGIC;
    rx_axis_tvalid_0 : OUT STD_LOGIC;
    rx_axis_tdata_0 : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
    rx_axis_tuser_0 : OUT STD_LOGIC_VECTOR(69 DOWNTO 0);
    ctl_rx_test_pattern_0 : IN STD_LOGIC;
    ctl_rx_enable_0 : IN STD_LOGIC;
    ctl_rx_delete_fcs_0 : IN STD_LOGIC;
    ctl_rx_ignore_fcs_0 : IN STD_LOGIC;
    ctl_rx_max_packet_len_0 : IN STD_LOGIC_VECTOR(14 DOWNTO 0);
    ctl_rx_min_packet_len_0 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    ctl_rx_custom_preamble_enable_0 : IN STD_LOGIC;
    ctl_rx_check_sfd_0 : IN STD_LOGIC;
    ctl_rx_check_preamble_0 : IN STD_LOGIC;
    ctl_rx_process_lfi_0 : IN STD_LOGIC;
    ctl_rx_force_resync_0 : IN STD_LOGIC;
    stat_rx_block_lock_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_framing_err_valid_0_0 : OUT STD_LOGIC;
    stat_rx_framing_err_0_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_1_0 : OUT STD_LOGIC;
    stat_rx_framing_err_1_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_2_0 : OUT STD_LOGIC;
    stat_rx_framing_err_2_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_3_0 : OUT STD_LOGIC;
    stat_rx_framing_err_3_0 : OUT STD_LOGIC;
    stat_rx_vl_demuxed_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_vl_number_0_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_1_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_2_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_3_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_synced_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_synced_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_len_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_repeat_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_misaligned_0 : OUT STD_LOGIC;
    stat_rx_aligned_err_0 : OUT STD_LOGIC;
    stat_rx_bip_err_0_0 : OUT STD_LOGIC;
    stat_rx_bip_err_1_0 : OUT STD_LOGIC;
    stat_rx_bip_err_2_0 : OUT STD_LOGIC;
    stat_rx_bip_err_3_0 : OUT STD_LOGIC;
    stat_rx_aligned_0 : OUT STD_LOGIC;
    stat_rx_hi_ber_0 : OUT STD_LOGIC;
    stat_rx_status_0 : OUT STD_LOGIC;
    stat_rx_bad_code_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_total_packets_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_total_good_packets_0 : OUT STD_LOGIC;
    stat_rx_total_bytes_0 : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    stat_rx_total_good_bytes_0 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_rx_packet_small_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_jabber_0 : OUT STD_LOGIC;
    stat_rx_packet_large_0 : OUT STD_LOGIC;
    stat_rx_oversize_0 : OUT STD_LOGIC;
    stat_rx_undersize_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_toolong_0 : OUT STD_LOGIC;
    stat_rx_fragment_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_64_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_65_127_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_128_255_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_256_511_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_512_1023_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1024_1518_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1519_1522_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1523_1548_bytes_0 : OUT STD_LOGIC;
    stat_rx_bad_fcs_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_bad_fcs_0 : OUT STD_LOGIC;
    stat_rx_stomped_fcs_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_1549_2047_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_2048_4095_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_4096_8191_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_8192_9215_bytes_0 : OUT STD_LOGIC;
    stat_rx_bad_preamble_0 : OUT STD_LOGIC;
    stat_rx_bad_sfd_0 : OUT STD_LOGIC;
    stat_rx_got_signal_os_0 : OUT STD_LOGIC;
    stat_rx_test_pattern_mismatch_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_truncated_0 : OUT STD_LOGIC;
    stat_rx_local_fault_0 : OUT STD_LOGIC;
    stat_rx_remote_fault_0 : OUT STD_LOGIC;
    stat_rx_internal_local_fault_0 : OUT STD_LOGIC;
    stat_rx_received_local_fault_0 : OUT STD_LOGIC;
    tx_reset_0 : IN STD_LOGIC;
    user_tx_reset_0 : OUT STD_LOGIC;
    tx_unfout_0 : OUT STD_LOGIC;
    tx_axis_tready_0 : OUT STD_LOGIC;
    tx_axis_tvalid_0 : IN STD_LOGIC;
    tx_axis_tdata_0 : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
    tx_axis_tuser_0 : IN STD_LOGIC_VECTOR(69 DOWNTO 0);
    stat_tx_total_packets_0 : OUT STD_LOGIC;
    stat_tx_total_bytes_0 : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
    stat_tx_total_good_packets_0 : OUT STD_LOGIC;
    stat_tx_total_good_bytes_0 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_tx_packet_64_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_65_127_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_128_255_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_256_511_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_512_1023_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1024_1518_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1519_1522_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1523_1548_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_small_0 : OUT STD_LOGIC;
    stat_tx_packet_large_0 : OUT STD_LOGIC;
    stat_tx_packet_1549_2047_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_2048_4095_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_4096_8191_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_8192_9215_bytes_0 : OUT STD_LOGIC;
    stat_tx_bad_fcs_0 : OUT STD_LOGIC;
    stat_tx_frame_error_0 : OUT STD_LOGIC;
    stat_tx_local_fault_0 : OUT STD_LOGIC;
    ctl_tx_test_pattern_0 : IN STD_LOGIC;
    ctl_tx_enable_0 : IN STD_LOGIC;
    ctl_tx_fcs_ins_enable_0 : IN STD_LOGIC;
    ctl_tx_ipg_value_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    ctl_tx_send_lfi_0 : IN STD_LOGIC;
    ctl_tx_send_rfi_0 : IN STD_LOGIC;
    ctl_tx_send_idle_0 : IN STD_LOGIC;
    ctl_tx_custom_preamble_enable_0 : IN STD_LOGIC;
    ctl_tx_ignore_fcs_0 : IN STD_LOGIC;
    gt_loopback_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    rx_core_clk_0 : IN STD_LOGIC
  );
END COMPONENT;


COMPONENT mac_40g_quad_132
  PORT (
    gt_rxp_in_0 : IN STD_LOGIC;
    gt_rxp_in_1 : IN STD_LOGIC;
    gt_rxp_in_2 : IN STD_LOGIC;
    gt_rxp_in_3 : IN STD_LOGIC;
    gt_rxn_in_0 : IN STD_LOGIC;
    gt_rxn_in_1 : IN STD_LOGIC;
    gt_rxn_in_2 : IN STD_LOGIC;
    gt_rxn_in_3 : IN STD_LOGIC;
    gt_txp_out_0 : OUT STD_LOGIC;
    gt_txp_out_1 : OUT STD_LOGIC;
    gt_txp_out_2 : OUT STD_LOGIC;
    gt_txp_out_3 : OUT STD_LOGIC;
    gt_txn_out_0 : OUT STD_LOGIC;
    gt_txn_out_1 : OUT STD_LOGIC;
    gt_txn_out_2 : OUT STD_LOGIC;
    gt_txn_out_3 : OUT STD_LOGIC;
    txoutclksel_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    rxoutclksel_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_dmonitorout_0 : OUT STD_LOGIC_VECTOR(67 DOWNTO 0);
    gt_eyescandataerror_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_eyescanreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_eyescantrigger_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_pcsrsvdin_0 : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
    gt_rxbufreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxbufstatus_0 : OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_rxcdrhold_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxcommadeten_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxdfeagchold_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxdfelpmreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxlatclk_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxlpmen_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpcsreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpmareset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpolarity_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbscntreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbserr_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbssel_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_rxrate_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_rxslide_in_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxstartofseq_0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    gt_txbufstatus_0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    gt_txdiffctrl_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gt_txinhibit_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txlatclk_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txmaincursor_0 : IN STD_LOGIC_VECTOR(27 DOWNTO 0);
    gt_txpcsreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpmareset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpolarity_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpostcursor_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gt_txprbsforceerr_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txprbssel_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_txprecursor_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gtwiz_reset_tx_datapath_0 : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    gtwiz_reset_rx_datapath_0 : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    rxrecclkout_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_common_drpclk : IN STD_LOGIC;
    gt_common_drpdo : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_common_drprdy : OUT STD_LOGIC;
    gt_common_drpen : IN STD_LOGIC;
    gt_common_drpwe : IN STD_LOGIC;
    gt_common_drpaddr : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_common_drpdi : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpclk_0 : IN STD_LOGIC;
    gt_ch_drpclk_1 : IN STD_LOGIC;
    gt_ch_drpclk_2 : IN STD_LOGIC;
    gt_ch_drpclk_3 : IN STD_LOGIC;
    gt_ch_drpdo_0 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_1 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_2 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_3 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drprdy_0 : OUT STD_LOGIC;
    gt_ch_drprdy_1 : OUT STD_LOGIC;
    gt_ch_drprdy_2 : OUT STD_LOGIC;
    gt_ch_drprdy_3 : OUT STD_LOGIC;
    gt_ch_drpen_0 : IN STD_LOGIC;
    gt_ch_drpen_1 : IN STD_LOGIC;
    gt_ch_drpen_2 : IN STD_LOGIC;
    gt_ch_drpen_3 : IN STD_LOGIC;
    gt_ch_drpwe_0 : IN STD_LOGIC;
    gt_ch_drpwe_1 : IN STD_LOGIC;
    gt_ch_drpwe_2 : IN STD_LOGIC;
    gt_ch_drpwe_3 : IN STD_LOGIC;
    gt_ch_drpaddr_0 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_1 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_2 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_3 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpdi_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_1 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_2 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_3 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    sys_reset : IN STD_LOGIC;
    dclk : IN STD_LOGIC;
    tx_clk_out_0 : OUT STD_LOGIC;
    rx_clk_out_0 : OUT STD_LOGIC;
    gt_refclk_p : IN STD_LOGIC;
    gt_refclk_n : IN STD_LOGIC;
    gt_refclk_out : OUT STD_LOGIC;
    gtpowergood_out_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    rx_reset_0 : IN STD_LOGIC;
    user_rx_reset_0 : OUT STD_LOGIC;
    rx_axis_tvalid_0 : OUT STD_LOGIC;
    rx_axis_tdata_0 : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
    rx_axis_tuser_0 : OUT STD_LOGIC_VECTOR(69 DOWNTO 0);
    ctl_rx_test_pattern_0 : IN STD_LOGIC;
    ctl_rx_enable_0 : IN STD_LOGIC;
    ctl_rx_delete_fcs_0 : IN STD_LOGIC;
    ctl_rx_ignore_fcs_0 : IN STD_LOGIC;
    ctl_rx_max_packet_len_0 : IN STD_LOGIC_VECTOR(14 DOWNTO 0);
    ctl_rx_min_packet_len_0 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    ctl_rx_custom_preamble_enable_0 : IN STD_LOGIC;
    ctl_rx_check_sfd_0 : IN STD_LOGIC;
    ctl_rx_check_preamble_0 : IN STD_LOGIC;
    ctl_rx_process_lfi_0 : IN STD_LOGIC;
    ctl_rx_force_resync_0 : IN STD_LOGIC;
    stat_rx_block_lock_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_framing_err_valid_0_0 : OUT STD_LOGIC;
    stat_rx_framing_err_0_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_1_0 : OUT STD_LOGIC;
    stat_rx_framing_err_1_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_2_0 : OUT STD_LOGIC;
    stat_rx_framing_err_2_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_3_0 : OUT STD_LOGIC;
    stat_rx_framing_err_3_0 : OUT STD_LOGIC;
    stat_rx_vl_demuxed_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_vl_number_0_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_1_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_2_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_3_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_synced_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_synced_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_len_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_repeat_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_misaligned_0 : OUT STD_LOGIC;
    stat_rx_aligned_err_0 : OUT STD_LOGIC;
    stat_rx_bip_err_0_0 : OUT STD_LOGIC;
    stat_rx_bip_err_1_0 : OUT STD_LOGIC;
    stat_rx_bip_err_2_0 : OUT STD_LOGIC;
    stat_rx_bip_err_3_0 : OUT STD_LOGIC;
    stat_rx_aligned_0 : OUT STD_LOGIC;
    stat_rx_hi_ber_0 : OUT STD_LOGIC;
    stat_rx_status_0 : OUT STD_LOGIC;
    stat_rx_bad_code_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_total_packets_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_total_good_packets_0 : OUT STD_LOGIC;
    stat_rx_total_bytes_0 : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    stat_rx_total_good_bytes_0 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_rx_packet_small_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_jabber_0 : OUT STD_LOGIC;
    stat_rx_packet_large_0 : OUT STD_LOGIC;
    stat_rx_oversize_0 : OUT STD_LOGIC;
    stat_rx_undersize_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_toolong_0 : OUT STD_LOGIC;
    stat_rx_fragment_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_64_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_65_127_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_128_255_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_256_511_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_512_1023_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1024_1518_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1519_1522_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1523_1548_bytes_0 : OUT STD_LOGIC;
    stat_rx_bad_fcs_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_bad_fcs_0 : OUT STD_LOGIC;
    stat_rx_stomped_fcs_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_1549_2047_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_2048_4095_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_4096_8191_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_8192_9215_bytes_0 : OUT STD_LOGIC;
    stat_rx_bad_preamble_0 : OUT STD_LOGIC;
    stat_rx_bad_sfd_0 : OUT STD_LOGIC;
    stat_rx_got_signal_os_0 : OUT STD_LOGIC;
    stat_rx_test_pattern_mismatch_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_truncated_0 : OUT STD_LOGIC;
    stat_rx_local_fault_0 : OUT STD_LOGIC;
    stat_rx_remote_fault_0 : OUT STD_LOGIC;
    stat_rx_internal_local_fault_0 : OUT STD_LOGIC;
    stat_rx_received_local_fault_0 : OUT STD_LOGIC;
    tx_reset_0 : IN STD_LOGIC;
    user_tx_reset_0 : OUT STD_LOGIC;
    tx_unfout_0 : OUT STD_LOGIC;
    tx_axis_tready_0 : OUT STD_LOGIC;
    tx_axis_tvalid_0 : IN STD_LOGIC;
    tx_axis_tdata_0 : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
    tx_axis_tuser_0 : IN STD_LOGIC_VECTOR(69 DOWNTO 0);
    stat_tx_total_packets_0 : OUT STD_LOGIC;
    stat_tx_total_bytes_0 : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
    stat_tx_total_good_packets_0 : OUT STD_LOGIC;
    stat_tx_total_good_bytes_0 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_tx_packet_64_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_65_127_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_128_255_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_256_511_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_512_1023_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1024_1518_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1519_1522_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1523_1548_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_small_0 : OUT STD_LOGIC;
    stat_tx_packet_large_0 : OUT STD_LOGIC;
    stat_tx_packet_1549_2047_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_2048_4095_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_4096_8191_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_8192_9215_bytes_0 : OUT STD_LOGIC;
    stat_tx_bad_fcs_0 : OUT STD_LOGIC;
    stat_tx_frame_error_0 : OUT STD_LOGIC;
    stat_tx_local_fault_0 : OUT STD_LOGIC;
    ctl_tx_test_pattern_0 : IN STD_LOGIC;
    ctl_tx_enable_0 : IN STD_LOGIC;
    ctl_tx_fcs_ins_enable_0 : IN STD_LOGIC;
    ctl_tx_ipg_value_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    ctl_tx_send_lfi_0 : IN STD_LOGIC;
    ctl_tx_send_rfi_0 : IN STD_LOGIC;
    ctl_tx_send_idle_0 : IN STD_LOGIC;
    ctl_tx_custom_preamble_enable_0 : IN STD_LOGIC;
    ctl_tx_ignore_fcs_0 : IN STD_LOGIC;
    gt_loopback_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    rx_core_clk_0 : IN STD_LOGIC
  );
END COMPONENT;


COMPONENT mac_40g_quad_134
  PORT (
    gt_rxp_in_0 : IN STD_LOGIC;
    gt_rxp_in_1 : IN STD_LOGIC;
    gt_rxp_in_2 : IN STD_LOGIC;
    gt_rxp_in_3 : IN STD_LOGIC;
    gt_rxn_in_0 : IN STD_LOGIC;
    gt_rxn_in_1 : IN STD_LOGIC;
    gt_rxn_in_2 : IN STD_LOGIC;
    gt_rxn_in_3 : IN STD_LOGIC;
    gt_txp_out_0 : OUT STD_LOGIC;
    gt_txp_out_1 : OUT STD_LOGIC;
    gt_txp_out_2 : OUT STD_LOGIC;
    gt_txp_out_3 : OUT STD_LOGIC;
    gt_txn_out_0 : OUT STD_LOGIC;
    gt_txn_out_1 : OUT STD_LOGIC;
    gt_txn_out_2 : OUT STD_LOGIC;
    gt_txn_out_3 : OUT STD_LOGIC;
    txoutclksel_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    rxoutclksel_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_dmonitorout_0 : OUT STD_LOGIC_VECTOR(67 DOWNTO 0);
    gt_eyescandataerror_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_eyescanreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_eyescantrigger_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_pcsrsvdin_0 : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
    gt_rxbufreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxbufstatus_0 : OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_rxcdrhold_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxcommadeten_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxdfeagchold_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxdfelpmreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxlatclk_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxlpmen_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpcsreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpmareset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpolarity_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbscntreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbserr_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbssel_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_rxrate_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_rxslide_in_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxstartofseq_0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    gt_txbufstatus_0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    gt_txdiffctrl_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gt_txinhibit_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txlatclk_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txmaincursor_0 : IN STD_LOGIC_VECTOR(27 DOWNTO 0);
    gt_txpcsreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpmareset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpolarity_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpostcursor_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gt_txprbsforceerr_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txprbssel_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_txprecursor_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gtwiz_reset_tx_datapath_0 : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    gtwiz_reset_rx_datapath_0 : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    rxrecclkout_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_common_drpclk : IN STD_LOGIC;
    gt_common_drpdo : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_common_drprdy : OUT STD_LOGIC;
    gt_common_drpen : IN STD_LOGIC;
    gt_common_drpwe : IN STD_LOGIC;
    gt_common_drpaddr : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_common_drpdi : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpclk_0 : IN STD_LOGIC;
    gt_ch_drpclk_1 : IN STD_LOGIC;
    gt_ch_drpclk_2 : IN STD_LOGIC;
    gt_ch_drpclk_3 : IN STD_LOGIC;
    gt_ch_drpdo_0 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_1 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_2 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_3 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drprdy_0 : OUT STD_LOGIC;
    gt_ch_drprdy_1 : OUT STD_LOGIC;
    gt_ch_drprdy_2 : OUT STD_LOGIC;
    gt_ch_drprdy_3 : OUT STD_LOGIC;
    gt_ch_drpen_0 : IN STD_LOGIC;
    gt_ch_drpen_1 : IN STD_LOGIC;
    gt_ch_drpen_2 : IN STD_LOGIC;
    gt_ch_drpen_3 : IN STD_LOGIC;
    gt_ch_drpwe_0 : IN STD_LOGIC;
    gt_ch_drpwe_1 : IN STD_LOGIC;
    gt_ch_drpwe_2 : IN STD_LOGIC;
    gt_ch_drpwe_3 : IN STD_LOGIC;
    gt_ch_drpaddr_0 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_1 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_2 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_3 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpdi_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_1 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_2 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_3 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    sys_reset : IN STD_LOGIC;
    dclk : IN STD_LOGIC;
    tx_clk_out_0 : OUT STD_LOGIC;
    rx_clk_out_0 : OUT STD_LOGIC;
    gt_refclk_p : IN STD_LOGIC;
    gt_refclk_n : IN STD_LOGIC;
    gt_refclk_out : OUT STD_LOGIC;
    gtpowergood_out_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    rx_reset_0 : IN STD_LOGIC;
    user_rx_reset_0 : OUT STD_LOGIC;
    rx_axis_tvalid_0 : OUT STD_LOGIC;
    rx_axis_tdata_0 : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
    rx_axis_tuser_0 : OUT STD_LOGIC_VECTOR(69 DOWNTO 0);
    ctl_rx_test_pattern_0 : IN STD_LOGIC;
    ctl_rx_enable_0 : IN STD_LOGIC;
    ctl_rx_delete_fcs_0 : IN STD_LOGIC;
    ctl_rx_ignore_fcs_0 : IN STD_LOGIC;
    ctl_rx_max_packet_len_0 : IN STD_LOGIC_VECTOR(14 DOWNTO 0);
    ctl_rx_min_packet_len_0 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    ctl_rx_custom_preamble_enable_0 : IN STD_LOGIC;
    ctl_rx_check_sfd_0 : IN STD_LOGIC;
    ctl_rx_check_preamble_0 : IN STD_LOGIC;
    ctl_rx_process_lfi_0 : IN STD_LOGIC;
    ctl_rx_force_resync_0 : IN STD_LOGIC;
    stat_rx_block_lock_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_framing_err_valid_0_0 : OUT STD_LOGIC;
    stat_rx_framing_err_0_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_1_0 : OUT STD_LOGIC;
    stat_rx_framing_err_1_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_2_0 : OUT STD_LOGIC;
    stat_rx_framing_err_2_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_3_0 : OUT STD_LOGIC;
    stat_rx_framing_err_3_0 : OUT STD_LOGIC;
    stat_rx_vl_demuxed_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_vl_number_0_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_1_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_2_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_3_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_synced_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_synced_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_len_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_repeat_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_misaligned_0 : OUT STD_LOGIC;
    stat_rx_aligned_err_0 : OUT STD_LOGIC;
    stat_rx_bip_err_0_0 : OUT STD_LOGIC;
    stat_rx_bip_err_1_0 : OUT STD_LOGIC;
    stat_rx_bip_err_2_0 : OUT STD_LOGIC;
    stat_rx_bip_err_3_0 : OUT STD_LOGIC;
    stat_rx_aligned_0 : OUT STD_LOGIC;
    stat_rx_hi_ber_0 : OUT STD_LOGIC;
    stat_rx_status_0 : OUT STD_LOGIC;
    stat_rx_bad_code_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_total_packets_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_total_good_packets_0 : OUT STD_LOGIC;
    stat_rx_total_bytes_0 : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    stat_rx_total_good_bytes_0 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_rx_packet_small_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_jabber_0 : OUT STD_LOGIC;
    stat_rx_packet_large_0 : OUT STD_LOGIC;
    stat_rx_oversize_0 : OUT STD_LOGIC;
    stat_rx_undersize_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_toolong_0 : OUT STD_LOGIC;
    stat_rx_fragment_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_64_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_65_127_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_128_255_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_256_511_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_512_1023_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1024_1518_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1519_1522_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1523_1548_bytes_0 : OUT STD_LOGIC;
    stat_rx_bad_fcs_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_bad_fcs_0 : OUT STD_LOGIC;
    stat_rx_stomped_fcs_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_1549_2047_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_2048_4095_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_4096_8191_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_8192_9215_bytes_0 : OUT STD_LOGIC;
    stat_rx_bad_preamble_0 : OUT STD_LOGIC;
    stat_rx_bad_sfd_0 : OUT STD_LOGIC;
    stat_rx_got_signal_os_0 : OUT STD_LOGIC;
    stat_rx_test_pattern_mismatch_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_truncated_0 : OUT STD_LOGIC;
    stat_rx_local_fault_0 : OUT STD_LOGIC;
    stat_rx_remote_fault_0 : OUT STD_LOGIC;
    stat_rx_internal_local_fault_0 : OUT STD_LOGIC;
    stat_rx_received_local_fault_0 : OUT STD_LOGIC;
    tx_reset_0 : IN STD_LOGIC;
    user_tx_reset_0 : OUT STD_LOGIC;
    tx_unfout_0 : OUT STD_LOGIC;
    tx_axis_tready_0 : OUT STD_LOGIC;
    tx_axis_tvalid_0 : IN STD_LOGIC;
    tx_axis_tdata_0 : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
    tx_axis_tuser_0 : IN STD_LOGIC_VECTOR(69 DOWNTO 0);
    stat_tx_total_packets_0 : OUT STD_LOGIC;
    stat_tx_total_bytes_0 : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
    stat_tx_total_good_packets_0 : OUT STD_LOGIC;
    stat_tx_total_good_bytes_0 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_tx_packet_64_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_65_127_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_128_255_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_256_511_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_512_1023_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1024_1518_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1519_1522_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1523_1548_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_small_0 : OUT STD_LOGIC;
    stat_tx_packet_large_0 : OUT STD_LOGIC;
    stat_tx_packet_1549_2047_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_2048_4095_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_4096_8191_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_8192_9215_bytes_0 : OUT STD_LOGIC;
    stat_tx_bad_fcs_0 : OUT STD_LOGIC;
    stat_tx_frame_error_0 : OUT STD_LOGIC;
    stat_tx_local_fault_0 : OUT STD_LOGIC;
    ctl_tx_test_pattern_0 : IN STD_LOGIC;
    ctl_tx_enable_0 : IN STD_LOGIC;
    ctl_tx_fcs_ins_enable_0 : IN STD_LOGIC;
    ctl_tx_ipg_value_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    ctl_tx_send_lfi_0 : IN STD_LOGIC;
    ctl_tx_send_rfi_0 : IN STD_LOGIC;
    ctl_tx_send_idle_0 : IN STD_LOGIC;
    ctl_tx_custom_preamble_enable_0 : IN STD_LOGIC;
    ctl_tx_ignore_fcs_0 : IN STD_LOGIC;
    gt_loopback_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    rx_core_clk_0 : IN STD_LOGIC
  );
END COMPONENT;

COMPONENT mac_40g_quad_135
  PORT (
    gt_rxp_in_0 : IN STD_LOGIC;
    gt_rxp_in_1 : IN STD_LOGIC;
    gt_rxp_in_2 : IN STD_LOGIC;
    gt_rxp_in_3 : IN STD_LOGIC;
    gt_rxn_in_0 : IN STD_LOGIC;
    gt_rxn_in_1 : IN STD_LOGIC;
    gt_rxn_in_2 : IN STD_LOGIC;
    gt_rxn_in_3 : IN STD_LOGIC;
    gt_txp_out_0 : OUT STD_LOGIC;
    gt_txp_out_1 : OUT STD_LOGIC;
    gt_txp_out_2 : OUT STD_LOGIC;
    gt_txp_out_3 : OUT STD_LOGIC;
    gt_txn_out_0 : OUT STD_LOGIC;
    gt_txn_out_1 : OUT STD_LOGIC;
    gt_txn_out_2 : OUT STD_LOGIC;
    gt_txn_out_3 : OUT STD_LOGIC;
    txoutclksel_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    rxoutclksel_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_dmonitorout_0 : OUT STD_LOGIC_VECTOR(67 DOWNTO 0);
    gt_eyescandataerror_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_eyescanreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_eyescantrigger_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_pcsrsvdin_0 : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
    gt_rxbufreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxbufstatus_0 : OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_rxcdrhold_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxcommadeten_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxdfeagchold_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxdfelpmreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxlatclk_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxlpmen_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpcsreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpmareset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxpolarity_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbscntreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbserr_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbssel_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_rxrate_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    gt_rxslide_in_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxstartofseq_0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    gt_txbufstatus_0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    gt_txdiffctrl_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gt_txinhibit_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txlatclk_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txmaincursor_0 : IN STD_LOGIC_VECTOR(27 DOWNTO 0);
    gt_txpcsreset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpmareset_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpolarity_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txpostcursor_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gt_txprbsforceerr_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txprbssel_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_txprecursor_0 : IN STD_LOGIC_VECTOR(19 DOWNTO 0);
    gtwiz_reset_tx_datapath_0 : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    gtwiz_reset_rx_datapath_0 : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    rxrecclkout_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_common_drpclk : IN STD_LOGIC;
    gt_common_drpdo : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_common_drprdy : OUT STD_LOGIC;
    gt_common_drpen : IN STD_LOGIC;
    gt_common_drpwe : IN STD_LOGIC;
    gt_common_drpaddr : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_common_drpdi : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpclk_0 : IN STD_LOGIC;
    gt_ch_drpclk_1 : IN STD_LOGIC;
    gt_ch_drpclk_2 : IN STD_LOGIC;
    gt_ch_drpclk_3 : IN STD_LOGIC;
    gt_ch_drpdo_0 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_1 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_2 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdo_3 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drprdy_0 : OUT STD_LOGIC;
    gt_ch_drprdy_1 : OUT STD_LOGIC;
    gt_ch_drprdy_2 : OUT STD_LOGIC;
    gt_ch_drprdy_3 : OUT STD_LOGIC;
    gt_ch_drpen_0 : IN STD_LOGIC;
    gt_ch_drpen_1 : IN STD_LOGIC;
    gt_ch_drpen_2 : IN STD_LOGIC;
    gt_ch_drpen_3 : IN STD_LOGIC;
    gt_ch_drpwe_0 : IN STD_LOGIC;
    gt_ch_drpwe_1 : IN STD_LOGIC;
    gt_ch_drpwe_2 : IN STD_LOGIC;
    gt_ch_drpwe_3 : IN STD_LOGIC;
    gt_ch_drpaddr_0 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_1 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_2 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpaddr_3 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_ch_drpdi_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_1 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_2 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_ch_drpdi_3 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    sys_reset : IN STD_LOGIC;
    dclk : IN STD_LOGIC;
    tx_clk_out_0 : OUT STD_LOGIC;
    rx_clk_out_0 : OUT STD_LOGIC;
    gt_refclk_p : IN STD_LOGIC;
    gt_refclk_n : IN STD_LOGIC;
    gt_refclk_out : OUT STD_LOGIC;
    gtpowergood_out_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    rx_reset_0 : IN STD_LOGIC;
    user_rx_reset_0 : OUT STD_LOGIC;
    rx_axis_tvalid_0 : OUT STD_LOGIC;
    rx_axis_tdata_0 : OUT STD_LOGIC_VECTOR(127 DOWNTO 0);
    rx_axis_tuser_0 : OUT STD_LOGIC_VECTOR(69 DOWNTO 0);
    ctl_rx_test_pattern_0 : IN STD_LOGIC;
    ctl_rx_enable_0 : IN STD_LOGIC;
    ctl_rx_delete_fcs_0 : IN STD_LOGIC;
    ctl_rx_ignore_fcs_0 : IN STD_LOGIC;
    ctl_rx_max_packet_len_0 : IN STD_LOGIC_VECTOR(14 DOWNTO 0);
    ctl_rx_min_packet_len_0 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    ctl_rx_custom_preamble_enable_0 : IN STD_LOGIC;
    ctl_rx_check_sfd_0 : IN STD_LOGIC;
    ctl_rx_check_preamble_0 : IN STD_LOGIC;
    ctl_rx_process_lfi_0 : IN STD_LOGIC;
    ctl_rx_force_resync_0 : IN STD_LOGIC;
    stat_rx_block_lock_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_framing_err_valid_0_0 : OUT STD_LOGIC;
    stat_rx_framing_err_0_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_1_0 : OUT STD_LOGIC;
    stat_rx_framing_err_1_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_2_0 : OUT STD_LOGIC;
    stat_rx_framing_err_2_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_3_0 : OUT STD_LOGIC;
    stat_rx_framing_err_3_0 : OUT STD_LOGIC;
    stat_rx_vl_demuxed_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_vl_number_0_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_1_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_2_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_vl_number_3_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_synced_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_synced_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_len_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_repeat_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_mf_err_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_misaligned_0 : OUT STD_LOGIC;
    stat_rx_aligned_err_0 : OUT STD_LOGIC;
    stat_rx_bip_err_0_0 : OUT STD_LOGIC;
    stat_rx_bip_err_1_0 : OUT STD_LOGIC;
    stat_rx_bip_err_2_0 : OUT STD_LOGIC;
    stat_rx_bip_err_3_0 : OUT STD_LOGIC;
    stat_rx_aligned_0 : OUT STD_LOGIC;
    stat_rx_hi_ber_0 : OUT STD_LOGIC;
    stat_rx_status_0 : OUT STD_LOGIC;
    stat_rx_bad_code_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_total_packets_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_total_good_packets_0 : OUT STD_LOGIC;
    stat_rx_total_bytes_0 : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    stat_rx_total_good_bytes_0 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_rx_packet_small_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_jabber_0 : OUT STD_LOGIC;
    stat_rx_packet_large_0 : OUT STD_LOGIC;
    stat_rx_oversize_0 : OUT STD_LOGIC;
    stat_rx_undersize_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_toolong_0 : OUT STD_LOGIC;
    stat_rx_fragment_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_64_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_65_127_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_128_255_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_256_511_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_512_1023_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1024_1518_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1519_1522_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1523_1548_bytes_0 : OUT STD_LOGIC;
    stat_rx_bad_fcs_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_bad_fcs_0 : OUT STD_LOGIC;
    stat_rx_stomped_fcs_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_packet_1549_2047_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_2048_4095_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_4096_8191_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_8192_9215_bytes_0 : OUT STD_LOGIC;
    stat_rx_bad_preamble_0 : OUT STD_LOGIC;
    stat_rx_bad_sfd_0 : OUT STD_LOGIC;
    stat_rx_got_signal_os_0 : OUT STD_LOGIC;
    stat_rx_test_pattern_mismatch_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_truncated_0 : OUT STD_LOGIC;
    stat_rx_local_fault_0 : OUT STD_LOGIC;
    stat_rx_remote_fault_0 : OUT STD_LOGIC;
    stat_rx_internal_local_fault_0 : OUT STD_LOGIC;
    stat_rx_received_local_fault_0 : OUT STD_LOGIC;
    tx_reset_0 : IN STD_LOGIC;
    user_tx_reset_0 : OUT STD_LOGIC;
    tx_unfout_0 : OUT STD_LOGIC;
    tx_axis_tready_0 : OUT STD_LOGIC;
    tx_axis_tvalid_0 : IN STD_LOGIC;
    tx_axis_tdata_0 : IN STD_LOGIC_VECTOR(127 DOWNTO 0);
    tx_axis_tuser_0 : IN STD_LOGIC_VECTOR(69 DOWNTO 0);
    stat_tx_total_packets_0 : OUT STD_LOGIC;
    stat_tx_total_bytes_0 : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
    stat_tx_total_good_packets_0 : OUT STD_LOGIC;
    stat_tx_total_good_bytes_0 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_tx_packet_64_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_65_127_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_128_255_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_256_511_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_512_1023_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1024_1518_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1519_1522_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1523_1548_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_small_0 : OUT STD_LOGIC;
    stat_tx_packet_large_0 : OUT STD_LOGIC;
    stat_tx_packet_1549_2047_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_2048_4095_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_4096_8191_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_8192_9215_bytes_0 : OUT STD_LOGIC;
    stat_tx_bad_fcs_0 : OUT STD_LOGIC;
    stat_tx_frame_error_0 : OUT STD_LOGIC;
    stat_tx_local_fault_0 : OUT STD_LOGIC;
    ctl_tx_test_pattern_0 : IN STD_LOGIC;
    ctl_tx_enable_0 : IN STD_LOGIC;
    ctl_tx_fcs_ins_enable_0 : IN STD_LOGIC;
    ctl_tx_ipg_value_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    ctl_tx_send_lfi_0 : IN STD_LOGIC;
    ctl_tx_send_rfi_0 : IN STD_LOGIC;
    ctl_tx_send_idle_0 : IN STD_LOGIC;
    ctl_tx_custom_preamble_enable_0 : IN STD_LOGIC;
    ctl_tx_ignore_fcs_0 : IN STD_LOGIC;
    gt_loopback_in_0 : IN STD_LOGIC_VECTOR(11 DOWNTO 0);
    rx_core_clk_0 : IN STD_LOGIC
  );
END COMPONENT;

END tech_mac_40g_component_pkg;

