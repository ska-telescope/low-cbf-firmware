LIBRARY IEEE, technology_lib;
USE IEEE.std_logic_1164.ALL;
USE technology_lib.technology_pkg.ALL;


PACKAGE tech_mac_10g_pkg IS

   TYPE t_locations_10g IS (
      SINGLE_10G_124_0, SINGLE_10G_120_3, SINGLE_10G_226_2);


END tech_mac_10g_pkg;

