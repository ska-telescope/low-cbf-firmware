-------------------------------------------------------------------------------
-- Title      : Visibility Definition Package
-- Project    : 
-------------------------------------------------------------------------------
-- File       : visibility_pkg.vhd
-- Author     : William Kamp  <william.kamp@aut.ac.nz>
-- Company    : High Performance Computing Research Lab, Auckland University of Technology
-- Created    : 2017-10-31
-- Last update: 2018-02-23
-- Platform   : 
-- Standard   : VHDL'2008
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Copyright (c) 2017 High Performance Computing Research Lab, Auckland University of Technology
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2017-10-31  1.0      will    Created
-- 2019-09-19  2.0p     nabel   Ported to Perentie (removed float_pkg and LTA data types)
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;

package visibility_pkg is

    type t_mta_data_frame is record
        baseline    : unsigned(19 downto 0);
        DVC         : unsigned(19 downto 0);
        TCI         : unsigned(39 downto 0);
        CCI         : unsigned(31 downto 0);
        pol_YY_real : signed(31 downto 0);
        pol_YY_imag : signed(31 downto 0);
        pol_YX_real : signed(31 downto 0);
        pol_YX_imag : signed(31 downto 0);
        pol_XY_real : signed(31 downto 0);
        pol_XY_imag : signed(31 downto 0);
        pol_XX_real : signed(31 downto 0);
        pol_XX_imag : signed(31 downto 0);
    end record t_mta_data_frame;

    type t_visibility_context is record
        tdm_lap_start : std_logic;
        tdm_lap       : unsigned(7 downto 0);
        channel       : unsigned(15 downto 0);
        timestamp     : unsigned(31 downto 0);
    end record t_visibility_context;

    --autogen start decl
 --------------------------------------------------
 -- Auto-generated code below. You should not edit.
 -- Generated Fri Feb 23 16:51:24 2018
 --------------------------------------------------
type t_mta_data_frame_a is array(natural range <>) of t_mta_data_frame;

constant T_MTA_DATA_FRAME_ZERO : t_mta_data_frame := (
	baseline => (others => '0'),
	DVC => (others => '0'),
	TCI => (others => '0'),
	CCI => (others => '0'),
	pol_YY_real => (others => '0'),
	pol_YY_imag => (others => '0'),
	pol_YX_real => (others => '0'),
	pol_YX_imag => (others => '0'),
	pol_XY_real => (others => '0'),
	pol_XY_imag => (others => '0'),
	pol_XX_real => (others => '0'),
	pol_XX_imag => (others => '0')
	);

constant T_MTA_DATA_FRAME_DONT_CARE : t_mta_data_frame := (
	baseline => (others => '-'),
	DVC => (others => '-'),
	TCI => (others => '-'),
	CCI => (others => '-'),
	pol_YY_real => (others => '-'),
	pol_YY_imag => (others => '-'),
	pol_YX_real => (others => '-'),
	pol_YX_imag => (others => '-'),
	pol_XY_real => (others => '-'),
	pol_XY_imag => (others => '-'),
	pol_XX_real => (others => '-'),
	pol_XX_imag => (others => '-')
	);

constant T_MTA_DATA_FRAME_SLV_WIDTH : natural := 368;

subtype t_mta_data_frame_slv is std_logic_vector(367 downto 0);
function to_slv (rec : t_mta_data_frame) return t_mta_data_frame_slv;

function from_slv (slv : std_logic_vector) return t_mta_data_frame;

type t_visibility_context_a is array(natural range <>) of t_visibility_context;

constant T_VISIBILITY_CONTEXT_ZERO : t_visibility_context := (
	tdm_lap_start => '0',
	tdm_lap => (others => '0'),
	channel => (others => '0'),
	timestamp => (others => '0')
	);

constant T_VISIBILITY_CONTEXT_DONT_CARE : t_visibility_context := (
	tdm_lap_start => '-',
	tdm_lap => (others => '-'),
	channel => (others => '-'),
	timestamp => (others => '-')
	);

constant T_VISIBILITY_CONTEXT_SLV_WIDTH : natural := 57;

subtype t_visibility_context_slv is std_logic_vector(56 downto 0);
function to_slv (rec : t_visibility_context) return t_visibility_context_slv;

function from_slv (slv : std_logic_vector) return t_visibility_context;

 ------------------------------------------------------
 -- End of Autogenerated code. You may add yours below.
 ------------------------------------------------------
    --autogen end decl

end package visibility_pkg;

package body visibility_pkg is

    --autogen start body
 --------------------------------------------------
 -- Auto-generated code below. You should not edit.
 -- Generated Fri Feb 23 16:51:24 2018
 --------------------------------------------------
function to_slv (rec : t_mta_data_frame) return t_mta_data_frame_slv is
    variable slv : std_logic_vector(367 downto 0);
begin
    slv(31 downto 0) := std_logic_vector(rec.pol_XX_imag);
    slv(63 downto 32) := std_logic_vector(rec.pol_XX_real);
    slv(95 downto 64) := std_logic_vector(rec.pol_XY_imag);
    slv(127 downto 96) := std_logic_vector(rec.pol_XY_real);
    slv(159 downto 128) := std_logic_vector(rec.pol_YX_imag);
    slv(191 downto 160) := std_logic_vector(rec.pol_YX_real);
    slv(223 downto 192) := std_logic_vector(rec.pol_YY_imag);
    slv(255 downto 224) := std_logic_vector(rec.pol_YY_real);
    slv(287 downto 256) := std_logic_vector(rec.CCI);
    slv(327 downto 288) := std_logic_vector(rec.TCI);
    slv(347 downto 328) := std_logic_vector(rec.DVC);
    slv(367 downto 348) := std_logic_vector(rec.baseline);
return slv;
end function to_slv;

function from_slv (slv : std_logic_vector) return t_mta_data_frame is
    variable rec : t_mta_data_frame;
begin
    rec.pol_XX_imag := signed(slv(31 downto 0));
    rec.pol_XX_real := signed(slv(63 downto 32));
    rec.pol_XY_imag := signed(slv(95 downto 64));
    rec.pol_XY_real := signed(slv(127 downto 96));
    rec.pol_YX_imag := signed(slv(159 downto 128));
    rec.pol_YX_real := signed(slv(191 downto 160));
    rec.pol_YY_imag := signed(slv(223 downto 192));
    rec.pol_YY_real := signed(slv(255 downto 224));
    rec.CCI := unsigned(slv(287 downto 256));
    rec.TCI := unsigned(slv(327 downto 288));
    rec.DVC := unsigned(slv(347 downto 328));
    rec.baseline := unsigned(slv(367 downto 348));
return rec;
end function from_slv;

function to_slv (rec : t_visibility_context) return t_visibility_context_slv is
    variable slv : std_logic_vector(56 downto 0);
begin
    slv(31 downto 0) := std_logic_vector(rec.timestamp);
    slv(47 downto 32) := std_logic_vector(rec.channel);
    slv(55 downto 48) := std_logic_vector(rec.tdm_lap);
    slv(56) := rec.tdm_lap_start;
return slv;
end function to_slv;

function from_slv (slv : std_logic_vector) return t_visibility_context is
    variable rec : t_visibility_context;
begin
    rec.timestamp := unsigned(slv(31 downto 0));
    rec.channel := unsigned(slv(47 downto 32));
    rec.tdm_lap := unsigned(slv(55 downto 48));
    rec.tdm_lap_start := slv(56);
return rec;
end function from_slv;

 ------------------------------------------------------
 -- End of Autogenerated code. You may add yours below.
 ------------------------------------------------------
    --autogen end body

end package body visibility_pkg;
