-------------------------------------------------------------------------------
--
-- File Name: ip_pkg.vhd
-- Contributing Authors: Andrew Brown
-- Type: RTL
-- Created: Wed Jun 13 16:40:00 2018
-- Template Rev: 1.0
--
-- Title: Gemini XH IP Library (ES FPGA)
--
-- Description: IP Library for Gemini XH (ES FPGA)
--
--
-- Compiler options:
--
--
-- Dependencies:
--
--
--
-------------------------------------------------------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

PACKAGE ip_pkg IS



END ip_pkg;
