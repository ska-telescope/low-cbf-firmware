----------------------------------------------------------------------------------
-- Company: CSIRO - CASS 
-- Engineer: David Humphrey
-- 
-- Create Date: 06.12.2018 09:59:02 
-- Module Name: PSTFBTop - Behavioral
-- Overview: 
--  low.CBF PST filterbank
--  Filterbank with 12 FIR taps, 256 point FFT, oversampled by a ratio of 4/3.
--  Designed for the low.CBF PST beamformer.
--  Processes 6 parallel signals, each with 8 bit complex data (8 bit real + 8 bit imaginary).
--  
-- Supporting Code:
--  The Matlab model should be in the directory ../matlab_model
--  Key files:
--   * ../matlab_model/run_PSTFB.m 
--       Generates input files for the simulation, runs the matlab model and compares with simulation output.
--   * ../matlab_model/get_rom_coefficients.m
--       Generates ROM data used in the firmware. ROMs are initialised using .coe files.
--       "PSTFIRTapsX.coe" : X runs from 1 to 12, contents of the 12 ROMS used to store the FIR filter taps.
--
--  Supporting VHDL 
--   * PSTFBtesttop.vhd 
--      Top level module that can be used to build this in a standalone version.
--   * PSTFB_tb.vhd
--      testbench, reads input data generated by the matlab code, and generates output data in text files for analysis by the matlab code. 
--
-- Structure:
--
--  File Structure
--  --------------
--  Outline of the structure shown below. Excludes most .xci files for DSPs, RAMs and ROMs.
--
--    PSTFBTop.vhd : This file, 6 complex inputs, 12 FIR filter taps, 256 point FFT, critically sampled
--        |
--        +-- PSTFBmem.vhd   : Input memory for the filterbank, 12 blocks of memory chained together, see "step 2. Filterbank memory" below.
--        +-- fb_DSP.vhd     : 12 TAP FIR filter, see "3. FIR filter" below.
--        +-- PSTFFTwrapper.vhd : 256 point FFT. see "4. 256 point FFT" below.
--                |
--                +-- fft256_16bit.xci : standard Xilinx 256 point FFT
--
--  Resource Use
--  ------------
--  Approximate resource usage is 
--   LUTs = 10320
--   DSPs = 216
--   Registers = 16474
--   BRAMs (36K) = 30
--
--  Power (estimate based on related measurement on the zcu111 board)
--   about 1 W static, 3.5 W dynamic.
--   
--  -----------------------------------------------------------------------------------------------
--  Description
--  -----------
--
-- 1. Controlling state machine
--   The oversampling requires that data be written and read from the memories in a particular pattern.
--   The state maching arranges this.
--
-- 2. Filterbank Memory
--   The filterbank memory consists of 11 blocks of memory chained together.
--   The read data from each memory is used both by the FIR filter and to write to the next memory in the chain.
--   The read and write addresses are staggered by one clock for each memory, implemented as a 12 sample delay line on
--   the address. This makes the timing easy to meet for the  memory address signals (which would otherwise be high-fanout signals)
--   and also enables use of the adders in the DSPs for the FIR filter.  
--
-- 3. FIR filter
--   The FIR filter uses 12 DSPs for each of the 12 simultaneous samples (6 channels * 2 (re+im)) that are read from the memory.
--   So the FIR filter uses (12 DSPS) * (6 simultaneous samples) * (2 (re+im)) = 144 DSPs.
--   The filter is implemented entirely in DSPs. The PCOUT port on the DSP is used to send the result of the multiplication
--   to the next DSP in the chain, where it is added using the adder in the DSP. This scheme requires that the inputs to the
--   12 DSPs are staggered to account for the pipeline stage on the PCOUT port. The staggering is done by controlling the address
--   to the memories as described above.
--
-- 4. 256 point FFT
--   Standard Xilinx FFT. Some messy logic at the front to account for the delay inserted by the "real-time" mode.
-- 
-- 5. Reorder memory
--   Data out of the FFT is in bit reversed order. It is stored in a double buffer in order from low to high frequencies,
--   and the central 216 fine channels are read out.
--
-- Reset behaviour
--  After a reset, the first "FRAMESTODROP" frames output is suppressed.
--  With "FRAMESTODROP" set to the default (15), the first output will be based entirely on valid input data
--  i.e. it is assumed that the first 11 input frames are initialisation data.
--  (Note that every 12 input frames generates 16 output frames due to the oversampling).  
----------------------------------------------------------------------------------
library IEEE, common_lib, filterbanks_lib;
use IEEE.STD_LOGIC_1164.ALL;
use common_lib.common_pkg.all;
use IEEE.NUMERIC_STD.ALL;

entity PSTFBTop is
    generic(
        METABITS : integer := 64;     -- Width in bits of the meta_i and meta_o ports.
        FRAMESTODROP : integer := 15  -- Number of output frames to drop after a reset (to account for initialisation of the filterbank)
    );
    port(
        -- clock, target is 380 MHz
        clk         : in std_logic;
        rst         : in std_logic;
        FIRTapUse_i : in std_logic;   -- FIR Taps are double buffered, choose which set of TAPs to use.
        -- Data input, common valid signal, expects packets of 64 samples. 
        -- Requires at least 2 clocks idle time between packets.
        -- Due to oversampling, also requires on average 86 clocks between packets - specifically, no more than 3 packets in 258 clocks. 
        data0_i : in t_slv_8_arr(1 downto 0);  -- 6 Inputs, each complex data, 8 bit real, 8 bit imaginary.
        data1_i : in t_slv_8_arr(1 downto 0);
        data2_i : in t_slv_8_arr(1 downto 0);
        data3_i : in t_slv_8_arr(1 downto 0);
        data4_i : in t_slv_8_arr(1 downto 0);
        data5_i : in t_slv_8_arr(1 downto 0);
        meta_i  : in std_logic_vector((METABITS-1) downto 0);  -- Sampled on the first cycle of every third packet of valid_i. 
        valid_i : in std_logic;
        -- Data out; bursts of 216 clocks for each channel.
        data0_o : out t_slv_16_arr(1 downto 0);   -- 6 outputs, real and imaginary parts in (0) and (1) respectively;
        data1_o : out t_slv_16_arr(1 downto 0);
        data2_o : out t_slv_16_arr(1 downto 0);
        data3_o : out t_slv_16_arr(1 downto 0);
        data4_o : out t_slv_16_arr(1 downto 0);
        data5_o : out t_slv_16_arr(1 downto 0);
        meta_o  : out std_logic_vector((METABITS-1) downto 0);
        valid_o : out std_logic;
        -- Writing FIR Taps
        FIRTapData_i   : in std_logic_vector(17 downto 0);  -- For register writes of the filtertaps.
        FIRTapData_o   : out std_logic_vector(17 downto 0); -- For register reads of the filtertaps. 3 cycle latency from FIRTapAddr_i
        FIRTapAddr_i   : in std_logic_vector(11 downto 0);   -- 256 * 12 filter taps = 3072 total.
        FIRTapWE_i     : in std_logic;
        FIRTapClk      : in std_logic;
        FIRTapSelect_i : in std_logic  -- FIR Taps are double buffered; This selects the buffer to access for registers. Choose which buffer to use with FIRTapUse_i
    );
end PSTFBTop;

architecture Behavioral of PSTFBTop is
    
    -- Reorder memory
    -- 3 BRAMs, simple dual port, 2 cycle read latency.
    -- Tcl:
    --  create_ip -name blk_mem_gen -vendor xilinx.com -library ip -version 8.4 -module_name PSTFBReorderMem -dir C:/projects/perentie/xilinx_test_projects/filterbank_ip
    --  set_property -dict [list CONFIG.Component_Name {PSTFBReorderMem} CONFIG.Memory_Type {Simple_Dual_Port_RAM} CONFIG.Assume_Synchronous_Clk {true} CONFIG.Write_Width_A {192} CONFIG.Write_Depth_A {512} CONFIG.Read_Width_A {192} CONFIG.Operating_Mode_A {NO_CHANGE} CONFIG.Enable_A {Always_Enabled} CONFIG.Write_Width_B {192} CONFIG.Read_Width_B {192} CONFIG.Operating_Mode_B {READ_FIRST} CONFIG.Enable_B {Always_Enabled} CONFIG.Register_PortA_Output_of_Memory_Primitives {false} CONFIG.Register_PortB_Output_of_Memory_Primitives {true} CONFIG.Fill_Remaining_Memory_Locations {true} CONFIG.Port_B_Clock {100} CONFIG.Port_B_Enable_Rate {100} CONFIG.Collision_Warnings {GENERATE_X_ONLY} CONFIG.Disable_Collision_Warnings {true} CONFIG.Disable_Out_of_Range_Warnings {true}] [get_ips PSTFBReorderMem]
    component PSTFBReorderMem
    port (
        clka  : in std_logic;
        wea   : in std_logic_vector(0 downto 0);
        addra : in std_logic_vector(8 downto 0);
        dina  : in std_logic_vector(191 downto 0);
        clkb  : in std_logic;
        addrb : in std_logic_vector(8 downto 0);
        doutb : out std_logic_vector(191 downto 0));
    end component;
    
    
    type rdFSM_type is (waitTrigger, run, waitDone);
    signal rdFSM : rdFSM_type;
    
    signal fbWrAddr : std_logic_vector(8 downto 0);
    signal validDel1 : std_logic;
    signal wrTriggerAddr : std_logic_vector(8 downto 0);
    signal rdTrigger : std_logic_vector(8 downto 0);
    signal rdTriggerValid : std_logic;
    
    signal fbRdAddr : std_logic_vector(8 downto 0);
    signal fbRdCount : std_logic_vector(7 downto 0);
    signal fbRdWrEn : std_logic;
    
    signal wrData96 : std_logic_vector(95 downto 0);
    signal fbmemRdData : t_slv_96_arr(11 downto 0);
    signal fbmemFIRTaps : t_slv_18_arr(11 downto 0);
    
    -- The first index in fbtype is for the number of filters = 12 (6 channels * 2[real+imaginary]).
    -- The second index is for the number of FIR taps.
    type fbtype is array(11 downto 0) of t_slv_8_arr(11 downto 0); 
    signal FBRdData : fbtype; 
    signal FIRDout : t_slv_16_arr(11 downto 0);
    signal fftIndex : t_slv_8_arr(5 downto 0);
    
    signal startAdv : std_logic_vector(31 downto 0);
    signal startFFT : std_logic := '0';
    
    signal fftRealOut : t_slv_16_arr(5 downto 0);
    signal fftImagOut : t_slv_16_arr(5 downto 0);
    signal fftvalidOut : std_logic_vector(5 downto 0) := "000000";
    

    signal reorderDout : std_logic_vector(191 downto 0);
    signal reorderWE : std_logic_vector(0 downto 0);
    signal reorderWrAddr : std_logic_vector(7 downto 0);
    signal reorderWrAddrFull : std_logic_vector(8 downto 0);
    signal reorderRdAddr, reorderRdAddrDel1 : std_logic_vector(7 downto 0);
    signal reorderRdAddrFull : std_logic_vector(8 downto 0);
    signal bufSelectWr, bufSelectRd : std_logic := '0';
    signal reorderDin : std_logic_vector(191 downto 0);
    signal rdRunning : std_logic := '0';
    signal rdRunningDel1, rdRunningDel2, rdRunningDel3 : std_logic := '0';
    signal validOutDel1 : std_logic := '0';
    signal bufSelectRdDel1, bufSelectRdDel2 : std_logic := '0';    
    
    signal metaDel0, metaDel1, metaDel2, metaDel3, metaDel4, metaDel5, metaDel6 : std_logic_vector(METABITS+16-1 downto 0);
    signal getMeta : std_logic;
    signal metaValid : std_logic;
    signal outputCount : std_logic_vector(15 downto 0);
    signal frameCountOut : std_logic_vector(15 downto 0);
    signal rdAddrFrameCount : std_logic_vector(3 downto 0);
    signal rotation : std_logic_vector(1 downto 0);
    signal metaDel2Count, metaDel3Count : std_logic_vector(7 downto 0) := (others => '0');
    
begin
    
    ------------------------------------------------------------------------------------
    -- 1. Controlling state machine
    -- ----------------------------   
    
    process(clk)
    begin
        if rising_edge(clk) then
        
            -- This is the write address to the first memory in the chain.
            -- It just counts up. The memory is 512 deep, so it wraps periodically. 
            if rst = '1' then
                fbWrAddr <= (others => '0');
            elsif valid_i = '1' then
                fbWrAddr <= std_logic_vector(unsigned(fbWrAddr) + 1);
            end if;
            validDel1 <= valid_i;
            
            -- Triggering of the read process. Oversampled so the read start address steps by 3/4 * 256 = 192 samples
            --  write 255 done   -> read 0-255
            --  write 447        -> read 192-447
            --  write 127        -> read 384-127
            --  write 319        -> read 64-319
            --  write 511        -> read 256-511
            --  write 191        -> read 448-191  <--- On reset, this triggers the first filterbank output. This is so that the output is aligned after the first 3072 samples have come in. 
            --  write 383        -> read 128-383
            --  write 63         -> read 320-63
            -- Then the pattern repeats:
            --  write 255        -> read 0-255    etc.
            -- 
            if rst = '1' then
                wrTriggerAddr <= "011000000";  -- 192
                rdTriggerValid <= '0';
                rdTrigger <= "000000000";
                outputCount <= "0000000000000001"; -- Count of the output frames to be generated.
            elsif (validDel1 = '1' and valid_i = '0' and fbWrAddr = wrTriggerAddr) then
                -- One clock after the last write.
                rdTrigger <= std_logic_vector(unsigned(wrTriggerAddr) - 256);
                rdTriggerValid <= '1';
                wrTriggerAddr <= std_logic_vector(unsigned(wrTriggerAddr) + 192);
                outputCount <= std_logic_vector(unsigned(outputCount) + 1);
            elsif rdFSM = waitTrigger then
                rdTriggerValid <= '0';
            end if;
            
            -- Meta data together with outputCount go into a delay line, which is sampled at the output to put the appropriate meta data with the output data.
            if rst = '1' then
                getMeta <= '1';
                metaValid <= '0';
            elsif valid_i = '1' and validDel1 = '0' and getMeta = '1' then
                metaDel0 <= outputCount & meta_i;
                metaValid <= '1';
                getMeta <= '0';
            elsif (validDel1 = '1' and valid_i = '0' and fbWrAddr = wrTriggerAddr) then
                -- falling edge of valid_i, for every third packet (of 64 samples) (i.e. once every 192 samples).
                getMeta <= '1';
                metaValid <= '0';
            else
                metaValid <= '0';
            end if;

            if metaValid = '1' then
                metaDel1 <= metaDel0;
            end if;
            if startAdv(0) = '1' then
                metaDel2 <= metaDel1;
                metaDel2Count <= "11111111";
            elsif metaDel2Count /= "00000000" then
                metaDel2Count <= std_logic_vector(unsigned(metaDel2Count) - 1);
            end if;
                 
            if metaDel2Count = "00000001" then
                metaDel3 <= metaDel2;
                metaDel3Count <= "11111111";
            elsif metaDel3Count /= "00000000" then
                metaDel3Count <= std_logic_vector(unsigned(metaDel3Count) - 1);
            end if;
            
            if metaDel3Count = "00000001" then
                metaDel4 <= metaDel3;
            end if;

            -- Simple FSM to control reading
            if rst = '1' then
               rdFSM <= waitTrigger;
            else
               case rdFSM is
                   when waitTrigger =>
                       fbRdCount <= "00000000";
                       if rdTriggerValid = '1' then
                           rdFSM <= run;
                           fbRdAddr <= rdTrigger;
                           fbRdWrEn <= '1';
                       else
                           fbRdWrEn <= '0';
                       end if;
                       
                   when run =>
                       if (unsigned(fbRdCount) = 255) then
                           rdFSM <= waitDone;
                       end if;
                       if (unsigned(fbRdCount) = 191) then
                           fbRdWrEn <= '0';
                       end if;
                       fbRdCount <= std_logic_vector(unsigned(fbRdCount) + 1);
                       fbRdAddr <= std_logic_vector(unsigned(fbRdAddr) + 1);
                       
                   when waitDone => -- Extra idle state ensures idle time between FFTs. 
                      rdFSM <= waitTrigger;
                      fbRdWrEn <= '0';
                       
                   when others =>
                       rdFSM <= waitTrigger;
               end case;
           end if;

        end if;
    end process;

    ------------------------------------------------------------------------------------
    -- 2. Input Memory
    -- ---------------
    
    wrData96 <= data5_i(1) & data5_i(0) & data4_i(1) & data4_i(0) & data3_i(1) & data3_i(0) & data2_i(1) & data2_i(0) & data1_i(1) & data1_i(0) & data0_i(1) & data0_i(0);

    cmem : entity filterbanks_lib.PSTFBMem
    generic map (
        TAPS => 12)  -- Note only partially parameterized; modification needed to support anything other than 12.
    port map (
        clk         => clk,
        FIRTapUse_i => FIRTapUse_i,   -- in std_logic; FIR Taps are double buffered, choose which set of TAPs to use.
        -- Write data for the start of the chain
        wrData_i    => wrData96,      -- in(95:0);
        wrAddr_i    => fbWrAddr,      -- in(8:0);
        wrEn_i      => valid_i,       -- in std_logic; should be a burst of 4096 clocks.
        -- Read data, comes out 2 clocks after the first write.
        rdData_o    => fbmemRdData,   -- out array96bit_type(TAPS-1 downto 0); -- 64 bits wide, 12 taps simultaneously; First sample is wr_data_i delayed by 1 clock.
        rdAddr_i    => fbRdAddr,      -- in(8:0);
        rdWrEn_i    => fbRdWrEn,      -- in std_logic;
        -- Read FIR Taps
        romAddr_i   => fbRdCount,     -- in(7:0);
        coef_o      => fbmemFIRTaps,  -- out array18bit_type(TAPS-1 downto 0); -- 18 bits per filter tap.
        -- Writing FIR Taps
        FIRTapData_i   => FIRTapData_i,   -- in(17:0);  -- For register writes of the filtertaps.
        FIRTapData_o   => FIRTapData_o,   -- out(17:0); -- For register reads of the filtertaps. 3 cycle latency from FIRTapAddr_i
        FIRTapAddr_i   => FIRTapAddr_i,   -- in(11:0);  -- 256 * 12 filter taps = 3072 total.
        FIRTapWE_i     => FIRTapWE_i,     -- in std_logic;
        FIRTapClk      => FIRTapClk,      -- in std_logic;
        FIRTapSelect_i => FIRTapSelect_i  -- in std_logic; FIR Taps are double buffered; this selects the buffer to access for registers. Choose which buffer to use with FIRTapUse_i
    );    

    
    -------------------------------------------------------------------------------------
    -- 3. FIR filter
    -- -------------
    -- 12 instances, 6 channels * (real + imaginary). Same filter taps used for all.
    -- PISA low.CBF processes simultaneously 2 (real+imaginary) * 3 (stations) * 2 (polarisations) = 12
    -- 
    
    CsampleGen : for j in 0 to 11 generate  -- 12 filters
        coefGen : for k in 0 to 11 generate  -- 12 taps
            FBRdData(j)(k) <= FBmemRdData(k)((j*8 + 7) downto (j*8));
        end generate;
    end generate;
    
    sampleGen : for j in 0 to 11 generate
            
        FIR : entity filterbanks_lib.fb_DSP
        generic map (
            TAPS => 12)  -- The module instantiates this number of DSPs
        port map (
            clk    => clk,
            data_i => FBRdData(j),  -- in array8bit_type(11 downto 0);
            coef_i => FBmemFIRTaps, -- in array18bit_type(11 downto 0);
            data_o => FIRDout(j)    -- out(15:0)
        );
    
    end generate;
    
    -------------------------------------------------------------------------------------
    -- 4. FFT
    -- -----------------
    -- 6 x 256 point FFTs.
    
    process(clk)
    begin
        if rising_edge(clk) then
            if (rdFSM = waitTrigger) and (rdTriggerValid = '1') then
                startAdv(0) <= '1';
            else
                startAdv(0) <= '0';
            end if;
            
            startAdv(31 downto 1) <= startAdv(30 downto 0);
            startFFT <= startAdv(14); -- Delay accounts for the delay through the FIR filter 
            
        end if;
    end process;
    
    
    fftgen : for j in 0 to 5 generate
        
        fft256 : entity filterbanks_lib.PSTFFTwrapper
        port map (
            clk  => clk,
            -- Input
            real_i  => FIRDout(j*2),     -- in(15:0); 16 bit real data
            imag_i  => FIRDout(j*2 + 1), -- in(15:0); 16 bit imaginary data
            start_i => startFFT,         -- in std_logic; pulse high; one clock in advance of the data 
            -- Output
            real_o  => fftRealOut(j), -- out(15:0);
            imag_o  => fftImagOut(j), -- out(15:0);
            index_o => fftIndex(j),   -- out(7:0);
            valid_o => fftvalidOut(j) -- out std_logic
        );
    
    end generate;
    
    -------------------------------------------------------------------------------------
    -- 5. Reorder the output from bit-reversed to the central 216 channels, low to high frequency.
    -- Uses a simple dual port BRAM double buffer.
      
    process(clk)
    begin
        if rising_edge(clk) then
        
            if (fftvalidOut(0) = '1' and (signed(fftIndex(0)) > -109) and (signed(fftIndex(0)) < 108)) then
                reorderWE(0) <= '1';
            else
                reorderWE(0) <= '0';
            end if;
            reorderWrAddr <= std_logic_vector(signed(fftIndex(0)) + 108);
            reorderDin <= fftImagOut(5) & fftRealOut(5) & fftImagOut(4) & fftRealOut(4) & fftImagOut(3) & fftRealOut(3) & fftImagOut(2) & fftRealOut(2) & fftImagOut(1) & fftRealOut(1) & fftImagOut(0) & fftRealOut(0);
            
            -- Falling edge of validOut triggers reading of the data from the memory
            validOutDel1 <= fftvalidOut(0);
            if fftvalidOut(0) = '0' and validOutDel1 = '1' then
                reorderRdAddr <= "00000000";
                bufSelectWr <= not bufSelectWr;
                bufSelectRd <= bufSelectWr;
                rdRunning <= '1';
            elsif rdRunning = '1' then
                reorderRdAddr <= std_logic_vector(unsigned(reorderRdAddr) + 1);
                -- read address runs from 0 to 215
                if unsigned(reorderRdAddr) = 215 then
                    rdRunning <= '0';
                end if;
            end if;
            rdRunningDel1 <= rdRunning;
            rdRunningDel2 <= rdRunningDel1;
            rdRunningDel3 <= rdRunningDel2;
            
            bufSelectRdDel1 <= bufSelectRd;
            bufSelectRdDel2 <= bufSelectRdDel1;
            
            reorderRdAddrDel1 <= reorderRdAddr;
            
        end if;
    end process;
    
    reorderWrAddrFull <= bufSelectWr & reorderWrAddr;
    reorderRdAddrFull <= bufSelectRd & reorderRdAddr;
    
    reorderRAM : PSTFBReorderMem
    port map (
        clka  => clk,
        wea   => reorderWE,         -- in std_logic_vector(0 downto 0);
        addra => reorderWrAddrFull, -- in(8:0);
        dina  => reorderDin,        -- in(191:0);
        clkb  => clk,
        addrb => reorderRdAddrFull, -- in(8:0);
        doutb => reorderDout        -- out(191:0)
    );

    rdAddrFrameCount <= reorderRdAddrDel1(1 downto 0) & frameCountOut(1 downto 0);

    process(clk)
    begin
        if rising_edge(clk) then

            if rdRunning = '1' and rdRunningDel1 = '0' then
                frameCountOut <= metaDel4((METABITS+15) downto METABITS);  -- frameCountOut aligns with rdRunningDel1 
            end if;
            
            -- DC will have a reorderRdAddr of 108 (decimal)
            case rdAddrFrameCount is
                when "0000" => rotation <= "00";  -- rotation aligns with rdRunningDel2
                when "0001" => rotation <= "00";
                when "0010" => rotation <= "00";
                when "0011" => rotation <= "00";
                when "0100" => rotation <= "00";
                when "0101" => rotation <= "01";
                when "0110" => rotation <= "10";
                when "0111" => rotation <= "11";
                when "1000" => rotation <= "00";
                when "1001" => rotation <= "10";
                when "1010" => rotation <= "00";
                when "1011" => rotation <= "10";
                when "1100" => rotation <= "00";
                when "1101" => rotation <= "11";
                when "1110" => rotation <= "10";
                when others => rotation <= "01";
            end case;
        
            if rotation = "00" then
                data0_o(0) <= reorderDout(15 downto 0);  -- dataX_o aligns with rdRunningDel3
                data0_o(1) <= reorderDout(31 downto 16);
                data1_o(0) <= reorderDout(47 downto 32);
                data1_o(1) <= reorderDout(63 downto 48);
                data2_o(0) <= reorderDout(79 downto 64);
                data2_o(1) <= reorderDout(95 downto 80);
                data3_o(0) <= reorderDout(111 downto 96);
                data3_o(1) <= reorderDout(127 downto 112);
                data4_o(0) <= reorderDout(143 downto 128);
                data4_o(1) <= reorderDout(159 downto 144);
                data5_o(0) <= reorderDout(175 downto 160);
                data5_o(1) <= reorderDout(191 downto 176);
            elsif rotation = "01" then  -- rotate +90 degrees; real -> imaginary, imaginary -> -real
                data0_o(0) <= std_logic_vector(-signed(reorderDout(31 downto 16)));
                data0_o(1) <= reorderDout(15 downto 0);
                data1_o(0) <= std_logic_vector(-signed(reorderDout(63 downto 48)));
                data1_o(1) <= reorderDout(47 downto 32);
                data2_o(0) <= std_logic_vector(-signed(reorderDout(95 downto 80)));
                data2_o(1) <= reorderDout(79 downto 64);
                data3_o(0) <= std_logic_vector(-signed(reorderDout(127 downto 112)));
                data3_o(1) <= reorderDout(111 downto 96);
                data4_o(0) <= std_logic_vector(-signed(reorderDout(159 downto 144)));
                data4_o(1) <= reorderDout(143 downto 128);
                data5_o(0) <= std_logic_vector(-signed(reorderDout(191 downto 176)));
                data5_o(1) <= reorderDout(175 downto 160);
            elsif rotation = "10" then -- rotation 180 degrees; real -> -real, imaginary -> -imaginary
                data0_o(0) <= std_logic_vector(-signed(reorderDout(15 downto 0)));
                data0_o(1) <= std_logic_vector(-signed(reorderDout(31 downto 16)));
                data1_o(0) <= std_logic_vector(-signed(reorderDout(47 downto 32)));
                data1_o(1) <= std_logic_vector(-signed(reorderDout(63 downto 48)));
                data2_o(0) <= std_logic_vector(-signed(reorderDout(79 downto 64)));
                data2_o(1) <= std_logic_vector(-signed(reorderDout(95 downto 80)));
                data3_o(0) <= std_logic_vector(-signed(reorderDout(111 downto 96)));
                data3_o(1) <= std_logic_vector(-signed(reorderDout(127 downto 112)));
                data4_o(0) <= std_logic_vector(-signed(reorderDout(143 downto 128)));
                data4_o(1) <= std_logic_vector(-signed(reorderDout(159 downto 144)));
                data5_o(0) <= std_logic_vector(-signed(reorderDout(175 downto 160)));
                data5_o(1) <= std_logic_vector(-signed(reorderDout(191 downto 176)));
            else  -- rotation = "11"; rotation 270 degrees; real -> -imaginary, imaginary -> real
                data0_o(0) <= reorderDout(31 downto 16);
                data0_o(1) <= std_logic_vector(-signed(reorderDout(15 downto 0)));
                data1_o(0) <= reorderDout(63 downto 48);
                data1_o(1) <= std_logic_vector(-signed(reorderDout(47 downto 32)));
                data2_o(0) <= reorderDout(95 downto 80);
                data2_o(1) <= std_logic_vector(-signed(reorderDout(79 downto 64)));
                data3_o(0) <= reorderDout(127 downto 112);
                data3_o(1) <= std_logic_vector(-signed(reorderDout(111 downto 96)));
                data4_o(0) <= reorderDout(159 downto 144);
                data4_o(1) <= std_logic_vector(-signed(reorderDout(143 downto 128)));
                data5_o(0) <= reorderDout(191 downto 176);
                data5_o(1) <= std_logic_vector(-signed(reorderDout(175 downto 160)));
            end if;
            
            if (unsigned(frameCountOut) > FRAMESTODROP) then
                valid_o <= rdRunningDel2;
            else
                valid_o <= '0';
            end if;
            
            if rdRunningDel2 = '1' and rdRunningDel3 = '0' then
                meta_o <= metaDel4((METABITS-1) downto 0);
            end if;
            
        end if;
    end process;
    
end Behavioral;
