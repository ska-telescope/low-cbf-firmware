LIBRARY IEEE, technology_lib;
USE IEEE.std_logic_1164.ALL;
USE technology_lib.technology_pkg.ALL;


PACKAGE tech_hbm_component_pkg IS

COMPONENT hbm_left_full
  PORT (
    HBM_REF_CLK_0 : IN STD_LOGIC;
    AXI_00_ACLK : IN STD_LOGIC;
    AXI_00_ARESET_N : IN STD_LOGIC;
    AXI_00_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_00_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_00_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_00_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_00_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_00_ARVALID : IN STD_LOGIC;
    AXI_00_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_00_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_00_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_00_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_00_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_00_AWVALID : IN STD_LOGIC;
    AXI_00_RREADY : IN STD_LOGIC;
    AXI_00_BREADY : IN STD_LOGIC;
    AXI_00_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_00_WLAST : IN STD_LOGIC;
    AXI_00_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_00_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_00_WVALID : IN STD_LOGIC;
    AXI_01_ACLK : IN STD_LOGIC;
    AXI_01_ARESET_N : IN STD_LOGIC;
    AXI_01_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_01_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_01_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_01_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_01_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_01_ARVALID : IN STD_LOGIC;
    AXI_01_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_01_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_01_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_01_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_01_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_01_AWVALID : IN STD_LOGIC;
    AXI_01_RREADY : IN STD_LOGIC;
    AXI_01_BREADY : IN STD_LOGIC;
    AXI_01_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_01_WLAST : IN STD_LOGIC;
    AXI_01_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_01_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_01_WVALID : IN STD_LOGIC;
    AXI_02_ACLK : IN STD_LOGIC;
    AXI_02_ARESET_N : IN STD_LOGIC;
    AXI_02_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_02_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_02_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_02_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_02_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_02_ARVALID : IN STD_LOGIC;
    AXI_02_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_02_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_02_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_02_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_02_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_02_AWVALID : IN STD_LOGIC;
    AXI_02_RREADY : IN STD_LOGIC;
    AXI_02_BREADY : IN STD_LOGIC;
    AXI_02_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_02_WLAST : IN STD_LOGIC;
    AXI_02_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_02_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_02_WVALID : IN STD_LOGIC;
    AXI_03_ACLK : IN STD_LOGIC;
    AXI_03_ARESET_N : IN STD_LOGIC;
    AXI_03_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_03_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_03_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_03_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_03_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_03_ARVALID : IN STD_LOGIC;
    AXI_03_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_03_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_03_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_03_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_03_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_03_AWVALID : IN STD_LOGIC;
    AXI_03_RREADY : IN STD_LOGIC;
    AXI_03_BREADY : IN STD_LOGIC;
    AXI_03_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_03_WLAST : IN STD_LOGIC;
    AXI_03_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_03_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_03_WVALID : IN STD_LOGIC;
    AXI_04_ACLK : IN STD_LOGIC;
    AXI_04_ARESET_N : IN STD_LOGIC;
    AXI_04_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_04_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_04_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_04_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_04_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_04_ARVALID : IN STD_LOGIC;
    AXI_04_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_04_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_04_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_04_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_04_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_04_AWVALID : IN STD_LOGIC;
    AXI_04_RREADY : IN STD_LOGIC;
    AXI_04_BREADY : IN STD_LOGIC;
    AXI_04_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_04_WLAST : IN STD_LOGIC;
    AXI_04_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_04_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_04_WVALID : IN STD_LOGIC;
    AXI_05_ACLK : IN STD_LOGIC;
    AXI_05_ARESET_N : IN STD_LOGIC;
    AXI_05_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_05_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_05_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_05_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_05_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_05_ARVALID : IN STD_LOGIC;
    AXI_05_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_05_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_05_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_05_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_05_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_05_AWVALID : IN STD_LOGIC;
    AXI_05_RREADY : IN STD_LOGIC;
    AXI_05_BREADY : IN STD_LOGIC;
    AXI_05_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_05_WLAST : IN STD_LOGIC;
    AXI_05_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_05_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_05_WVALID : IN STD_LOGIC;
    AXI_06_ACLK : IN STD_LOGIC;
    AXI_06_ARESET_N : IN STD_LOGIC;
    AXI_06_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_06_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_06_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_06_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_06_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_06_ARVALID : IN STD_LOGIC;
    AXI_06_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_06_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_06_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_06_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_06_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_06_AWVALID : IN STD_LOGIC;
    AXI_06_RREADY : IN STD_LOGIC;
    AXI_06_BREADY : IN STD_LOGIC;
    AXI_06_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_06_WLAST : IN STD_LOGIC;
    AXI_06_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_06_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_06_WVALID : IN STD_LOGIC;
    AXI_07_ACLK : IN STD_LOGIC;
    AXI_07_ARESET_N : IN STD_LOGIC;
    AXI_07_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_07_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_07_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_07_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_07_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_07_ARVALID : IN STD_LOGIC;
    AXI_07_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_07_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_07_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_07_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_07_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_07_AWVALID : IN STD_LOGIC;
    AXI_07_RREADY : IN STD_LOGIC;
    AXI_07_BREADY : IN STD_LOGIC;
    AXI_07_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_07_WLAST : IN STD_LOGIC;
    AXI_07_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_07_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_07_WVALID : IN STD_LOGIC;
    AXI_08_ACLK : IN STD_LOGIC;
    AXI_08_ARESET_N : IN STD_LOGIC;
    AXI_08_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_08_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_08_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_08_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_08_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_08_ARVALID : IN STD_LOGIC;
    AXI_08_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_08_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_08_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_08_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_08_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_08_AWVALID : IN STD_LOGIC;
    AXI_08_RREADY : IN STD_LOGIC;
    AXI_08_BREADY : IN STD_LOGIC;
    AXI_08_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_08_WLAST : IN STD_LOGIC;
    AXI_08_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_08_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_08_WVALID : IN STD_LOGIC;
    AXI_09_ACLK : IN STD_LOGIC;
    AXI_09_ARESET_N : IN STD_LOGIC;
    AXI_09_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_09_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_09_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_09_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_09_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_09_ARVALID : IN STD_LOGIC;
    AXI_09_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_09_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_09_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_09_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_09_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_09_AWVALID : IN STD_LOGIC;
    AXI_09_RREADY : IN STD_LOGIC;
    AXI_09_BREADY : IN STD_LOGIC;
    AXI_09_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_09_WLAST : IN STD_LOGIC;
    AXI_09_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_09_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_09_WVALID : IN STD_LOGIC;
    AXI_10_ACLK : IN STD_LOGIC;
    AXI_10_ARESET_N : IN STD_LOGIC;
    AXI_10_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_10_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_10_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_10_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_10_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_10_ARVALID : IN STD_LOGIC;
    AXI_10_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_10_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_10_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_10_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_10_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_10_AWVALID : IN STD_LOGIC;
    AXI_10_RREADY : IN STD_LOGIC;
    AXI_10_BREADY : IN STD_LOGIC;
    AXI_10_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_10_WLAST : IN STD_LOGIC;
    AXI_10_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_10_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_10_WVALID : IN STD_LOGIC;
    AXI_11_ACLK : IN STD_LOGIC;
    AXI_11_ARESET_N : IN STD_LOGIC;
    AXI_11_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_11_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_11_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_11_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_11_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_11_ARVALID : IN STD_LOGIC;
    AXI_11_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_11_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_11_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_11_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_11_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_11_AWVALID : IN STD_LOGIC;
    AXI_11_RREADY : IN STD_LOGIC;
    AXI_11_BREADY : IN STD_LOGIC;
    AXI_11_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_11_WLAST : IN STD_LOGIC;
    AXI_11_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_11_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_11_WVALID : IN STD_LOGIC;
    AXI_12_ACLK : IN STD_LOGIC;
    AXI_12_ARESET_N : IN STD_LOGIC;
    AXI_12_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_12_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_12_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_12_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_12_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_12_ARVALID : IN STD_LOGIC;
    AXI_12_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_12_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_12_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_12_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_12_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_12_AWVALID : IN STD_LOGIC;
    AXI_12_RREADY : IN STD_LOGIC;
    AXI_12_BREADY : IN STD_LOGIC;
    AXI_12_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_12_WLAST : IN STD_LOGIC;
    AXI_12_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_12_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_12_WVALID : IN STD_LOGIC;
    AXI_13_ACLK : IN STD_LOGIC;
    AXI_13_ARESET_N : IN STD_LOGIC;
    AXI_13_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_13_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_13_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_13_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_13_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_13_ARVALID : IN STD_LOGIC;
    AXI_13_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_13_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_13_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_13_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_13_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_13_AWVALID : IN STD_LOGIC;
    AXI_13_RREADY : IN STD_LOGIC;
    AXI_13_BREADY : IN STD_LOGIC;
    AXI_13_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_13_WLAST : IN STD_LOGIC;
    AXI_13_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_13_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_13_WVALID : IN STD_LOGIC;
    AXI_14_ACLK : IN STD_LOGIC;
    AXI_14_ARESET_N : IN STD_LOGIC;
    AXI_14_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_14_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_14_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_14_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_14_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_14_ARVALID : IN STD_LOGIC;
    AXI_14_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_14_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_14_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_14_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_14_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_14_AWVALID : IN STD_LOGIC;
    AXI_14_RREADY : IN STD_LOGIC;
    AXI_14_BREADY : IN STD_LOGIC;
    AXI_14_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_14_WLAST : IN STD_LOGIC;
    AXI_14_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_14_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_14_WVALID : IN STD_LOGIC;
    AXI_15_ACLK : IN STD_LOGIC;
    AXI_15_ARESET_N : IN STD_LOGIC;
    AXI_15_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_15_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_15_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_15_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_15_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_15_ARVALID : IN STD_LOGIC;
    AXI_15_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_15_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_15_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_15_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_15_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_15_AWVALID : IN STD_LOGIC;
    AXI_15_RREADY : IN STD_LOGIC;
    AXI_15_BREADY : IN STD_LOGIC;
    AXI_15_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_15_WLAST : IN STD_LOGIC;
    AXI_15_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_15_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_15_WVALID : IN STD_LOGIC;
    APB_0_PWDATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    APB_0_PADDR : IN STD_LOGIC_VECTOR(21 DOWNTO 0);
    APB_0_PCLK : IN STD_LOGIC;
    APB_0_PENABLE : IN STD_LOGIC;
    APB_0_PRESET_N : IN STD_LOGIC;
    APB_0_PSEL : IN STD_LOGIC;
    APB_0_PWRITE : IN STD_LOGIC;
    AXI_00_ARREADY : OUT STD_LOGIC;
    AXI_00_AWREADY : OUT STD_LOGIC;
    AXI_00_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_00_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_00_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_00_RLAST : OUT STD_LOGIC;
    AXI_00_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_00_RVALID : OUT STD_LOGIC;
    AXI_00_WREADY : OUT STD_LOGIC;
    AXI_00_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_00_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_00_BVALID : OUT STD_LOGIC;
    AXI_01_ARREADY : OUT STD_LOGIC;
    AXI_01_AWREADY : OUT STD_LOGIC;
    AXI_01_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_01_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_01_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_01_RLAST : OUT STD_LOGIC;
    AXI_01_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_01_RVALID : OUT STD_LOGIC;
    AXI_01_WREADY : OUT STD_LOGIC;
    AXI_01_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_01_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_01_BVALID : OUT STD_LOGIC;
    AXI_02_ARREADY : OUT STD_LOGIC;
    AXI_02_AWREADY : OUT STD_LOGIC;
    AXI_02_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_02_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_02_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_02_RLAST : OUT STD_LOGIC;
    AXI_02_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_02_RVALID : OUT STD_LOGIC;
    AXI_02_WREADY : OUT STD_LOGIC;
    AXI_02_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_02_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_02_BVALID : OUT STD_LOGIC;
    AXI_03_ARREADY : OUT STD_LOGIC;
    AXI_03_AWREADY : OUT STD_LOGIC;
    AXI_03_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_03_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_03_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_03_RLAST : OUT STD_LOGIC;
    AXI_03_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_03_RVALID : OUT STD_LOGIC;
    AXI_03_WREADY : OUT STD_LOGIC;
    AXI_03_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_03_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_03_BVALID : OUT STD_LOGIC;
    AXI_04_ARREADY : OUT STD_LOGIC;
    AXI_04_AWREADY : OUT STD_LOGIC;
    AXI_04_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_04_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_04_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_04_RLAST : OUT STD_LOGIC;
    AXI_04_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_04_RVALID : OUT STD_LOGIC;
    AXI_04_WREADY : OUT STD_LOGIC;
    AXI_04_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_04_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_04_BVALID : OUT STD_LOGIC;
    AXI_05_ARREADY : OUT STD_LOGIC;
    AXI_05_AWREADY : OUT STD_LOGIC;
    AXI_05_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_05_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_05_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_05_RLAST : OUT STD_LOGIC;
    AXI_05_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_05_RVALID : OUT STD_LOGIC;
    AXI_05_WREADY : OUT STD_LOGIC;
    AXI_05_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_05_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_05_BVALID : OUT STD_LOGIC;
    AXI_06_ARREADY : OUT STD_LOGIC;
    AXI_06_AWREADY : OUT STD_LOGIC;
    AXI_06_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_06_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_06_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_06_RLAST : OUT STD_LOGIC;
    AXI_06_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_06_RVALID : OUT STD_LOGIC;
    AXI_06_WREADY : OUT STD_LOGIC;
    AXI_06_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_06_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_06_BVALID : OUT STD_LOGIC;
    AXI_07_ARREADY : OUT STD_LOGIC;
    AXI_07_AWREADY : OUT STD_LOGIC;
    AXI_07_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_07_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_07_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_07_RLAST : OUT STD_LOGIC;
    AXI_07_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_07_RVALID : OUT STD_LOGIC;
    AXI_07_WREADY : OUT STD_LOGIC;
    AXI_07_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_07_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_07_BVALID : OUT STD_LOGIC;
    AXI_08_ARREADY : OUT STD_LOGIC;
    AXI_08_AWREADY : OUT STD_LOGIC;
    AXI_08_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_08_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_08_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_08_RLAST : OUT STD_LOGIC;
    AXI_08_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_08_RVALID : OUT STD_LOGIC;
    AXI_08_WREADY : OUT STD_LOGIC;
    AXI_08_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_08_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_08_BVALID : OUT STD_LOGIC;
    AXI_09_ARREADY : OUT STD_LOGIC;
    AXI_09_AWREADY : OUT STD_LOGIC;
    AXI_09_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_09_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_09_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_09_RLAST : OUT STD_LOGIC;
    AXI_09_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_09_RVALID : OUT STD_LOGIC;
    AXI_09_WREADY : OUT STD_LOGIC;
    AXI_09_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_09_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_09_BVALID : OUT STD_LOGIC;
    AXI_10_ARREADY : OUT STD_LOGIC;
    AXI_10_AWREADY : OUT STD_LOGIC;
    AXI_10_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_10_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_10_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_10_RLAST : OUT STD_LOGIC;
    AXI_10_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_10_RVALID : OUT STD_LOGIC;
    AXI_10_WREADY : OUT STD_LOGIC;
    AXI_10_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_10_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_10_BVALID : OUT STD_LOGIC;
    AXI_11_ARREADY : OUT STD_LOGIC;
    AXI_11_AWREADY : OUT STD_LOGIC;
    AXI_11_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_11_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_11_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_11_RLAST : OUT STD_LOGIC;
    AXI_11_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_11_RVALID : OUT STD_LOGIC;
    AXI_11_WREADY : OUT STD_LOGIC;
    AXI_11_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_11_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_11_BVALID : OUT STD_LOGIC;
    AXI_12_ARREADY : OUT STD_LOGIC;
    AXI_12_AWREADY : OUT STD_LOGIC;
    AXI_12_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_12_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_12_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_12_RLAST : OUT STD_LOGIC;
    AXI_12_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_12_RVALID : OUT STD_LOGIC;
    AXI_12_WREADY : OUT STD_LOGIC;
    AXI_12_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_12_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_12_BVALID : OUT STD_LOGIC;
    AXI_13_ARREADY : OUT STD_LOGIC;
    AXI_13_AWREADY : OUT STD_LOGIC;
    AXI_13_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_13_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_13_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_13_RLAST : OUT STD_LOGIC;
    AXI_13_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_13_RVALID : OUT STD_LOGIC;
    AXI_13_WREADY : OUT STD_LOGIC;
    AXI_13_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_13_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_13_BVALID : OUT STD_LOGIC;
    AXI_14_ARREADY : OUT STD_LOGIC;
    AXI_14_AWREADY : OUT STD_LOGIC;
    AXI_14_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_14_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_14_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_14_RLAST : OUT STD_LOGIC;
    AXI_14_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_14_RVALID : OUT STD_LOGIC;
    AXI_14_WREADY : OUT STD_LOGIC;
    AXI_14_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_14_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_14_BVALID : OUT STD_LOGIC;
    AXI_15_ARREADY : OUT STD_LOGIC;
    AXI_15_AWREADY : OUT STD_LOGIC;
    AXI_15_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_15_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_15_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_15_RLAST : OUT STD_LOGIC;
    AXI_15_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_15_RVALID : OUT STD_LOGIC;
    AXI_15_WREADY : OUT STD_LOGIC;
    AXI_15_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_15_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_15_BVALID : OUT STD_LOGIC;
    APB_0_PRDATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    APB_0_PREADY : OUT STD_LOGIC;
    APB_0_PSLVERR : OUT STD_LOGIC;
    apb_complete_0 : OUT STD_LOGIC;
    DRAM_0_STAT_CATTRIP : OUT STD_LOGIC;
    DRAM_0_STAT_TEMP : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
  );
END COMPONENT;


COMPONENT hbm_right_individual
  PORT (
    HBM_REF_CLK_0 : IN STD_LOGIC;
    AXI_00_ACLK : IN STD_LOGIC;
    AXI_00_ARESET_N : IN STD_LOGIC;
    AXI_00_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_00_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_00_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_00_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_00_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_00_ARVALID : IN STD_LOGIC;
    AXI_00_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_00_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_00_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_00_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_00_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_00_AWVALID : IN STD_LOGIC;
    AXI_00_RREADY : IN STD_LOGIC;
    AXI_00_BREADY : IN STD_LOGIC;
    AXI_00_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_00_WLAST : IN STD_LOGIC;
    AXI_00_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_00_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_00_WVALID : IN STD_LOGIC;
    AXI_01_ACLK : IN STD_LOGIC;
    AXI_01_ARESET_N : IN STD_LOGIC;
    AXI_01_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_01_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_01_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_01_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_01_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_01_ARVALID : IN STD_LOGIC;
    AXI_01_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_01_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_01_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_01_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_01_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_01_AWVALID : IN STD_LOGIC;
    AXI_01_RREADY : IN STD_LOGIC;
    AXI_01_BREADY : IN STD_LOGIC;
    AXI_01_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_01_WLAST : IN STD_LOGIC;
    AXI_01_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_01_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_01_WVALID : IN STD_LOGIC;
    AXI_02_ACLK : IN STD_LOGIC;
    AXI_02_ARESET_N : IN STD_LOGIC;
    AXI_02_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_02_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_02_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_02_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_02_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_02_ARVALID : IN STD_LOGIC;
    AXI_02_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_02_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_02_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_02_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_02_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_02_AWVALID : IN STD_LOGIC;
    AXI_02_RREADY : IN STD_LOGIC;
    AXI_02_BREADY : IN STD_LOGIC;
    AXI_02_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_02_WLAST : IN STD_LOGIC;
    AXI_02_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_02_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_02_WVALID : IN STD_LOGIC;
    AXI_03_ACLK : IN STD_LOGIC;
    AXI_03_ARESET_N : IN STD_LOGIC;
    AXI_03_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_03_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_03_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_03_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_03_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_03_ARVALID : IN STD_LOGIC;
    AXI_03_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_03_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_03_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_03_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_03_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_03_AWVALID : IN STD_LOGIC;
    AXI_03_RREADY : IN STD_LOGIC;
    AXI_03_BREADY : IN STD_LOGIC;
    AXI_03_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_03_WLAST : IN STD_LOGIC;
    AXI_03_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_03_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_03_WVALID : IN STD_LOGIC;
    AXI_04_ACLK : IN STD_LOGIC;
    AXI_04_ARESET_N : IN STD_LOGIC;
    AXI_04_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_04_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_04_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_04_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_04_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_04_ARVALID : IN STD_LOGIC;
    AXI_04_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_04_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_04_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_04_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_04_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_04_AWVALID : IN STD_LOGIC;
    AXI_04_RREADY : IN STD_LOGIC;
    AXI_04_BREADY : IN STD_LOGIC;
    AXI_04_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_04_WLAST : IN STD_LOGIC;
    AXI_04_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_04_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_04_WVALID : IN STD_LOGIC;
    AXI_05_ACLK : IN STD_LOGIC;
    AXI_05_ARESET_N : IN STD_LOGIC;
    AXI_05_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_05_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_05_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_05_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_05_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_05_ARVALID : IN STD_LOGIC;
    AXI_05_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_05_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_05_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_05_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_05_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_05_AWVALID : IN STD_LOGIC;
    AXI_05_RREADY : IN STD_LOGIC;
    AXI_05_BREADY : IN STD_LOGIC;
    AXI_05_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_05_WLAST : IN STD_LOGIC;
    AXI_05_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_05_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_05_WVALID : IN STD_LOGIC;
    AXI_06_ACLK : IN STD_LOGIC;
    AXI_06_ARESET_N : IN STD_LOGIC;
    AXI_06_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_06_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_06_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_06_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_06_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_06_ARVALID : IN STD_LOGIC;
    AXI_06_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_06_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_06_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_06_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_06_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_06_AWVALID : IN STD_LOGIC;
    AXI_06_RREADY : IN STD_LOGIC;
    AXI_06_BREADY : IN STD_LOGIC;
    AXI_06_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_06_WLAST : IN STD_LOGIC;
    AXI_06_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_06_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_06_WVALID : IN STD_LOGIC;
    AXI_07_ACLK : IN STD_LOGIC;
    AXI_07_ARESET_N : IN STD_LOGIC;
    AXI_07_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_07_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_07_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_07_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_07_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_07_ARVALID : IN STD_LOGIC;
    AXI_07_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_07_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_07_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_07_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_07_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_07_AWVALID : IN STD_LOGIC;
    AXI_07_RREADY : IN STD_LOGIC;
    AXI_07_BREADY : IN STD_LOGIC;
    AXI_07_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_07_WLAST : IN STD_LOGIC;
    AXI_07_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_07_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_07_WVALID : IN STD_LOGIC;
    AXI_08_ACLK : IN STD_LOGIC;
    AXI_08_ARESET_N : IN STD_LOGIC;
    AXI_08_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_08_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_08_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_08_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_08_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_08_ARVALID : IN STD_LOGIC;
    AXI_08_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_08_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_08_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_08_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_08_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_08_AWVALID : IN STD_LOGIC;
    AXI_08_RREADY : IN STD_LOGIC;
    AXI_08_BREADY : IN STD_LOGIC;
    AXI_08_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_08_WLAST : IN STD_LOGIC;
    AXI_08_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_08_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_08_WVALID : IN STD_LOGIC;
    AXI_09_ACLK : IN STD_LOGIC;
    AXI_09_ARESET_N : IN STD_LOGIC;
    AXI_09_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_09_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_09_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_09_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_09_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_09_ARVALID : IN STD_LOGIC;
    AXI_09_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_09_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_09_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_09_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_09_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_09_AWVALID : IN STD_LOGIC;
    AXI_09_RREADY : IN STD_LOGIC;
    AXI_09_BREADY : IN STD_LOGIC;
    AXI_09_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_09_WLAST : IN STD_LOGIC;
    AXI_09_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_09_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_09_WVALID : IN STD_LOGIC;
    AXI_10_ACLK : IN STD_LOGIC;
    AXI_10_ARESET_N : IN STD_LOGIC;
    AXI_10_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_10_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_10_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_10_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_10_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_10_ARVALID : IN STD_LOGIC;
    AXI_10_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_10_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_10_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_10_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_10_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_10_AWVALID : IN STD_LOGIC;
    AXI_10_RREADY : IN STD_LOGIC;
    AXI_10_BREADY : IN STD_LOGIC;
    AXI_10_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_10_WLAST : IN STD_LOGIC;
    AXI_10_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_10_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_10_WVALID : IN STD_LOGIC;
    AXI_11_ACLK : IN STD_LOGIC;
    AXI_11_ARESET_N : IN STD_LOGIC;
    AXI_11_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_11_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_11_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_11_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_11_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_11_ARVALID : IN STD_LOGIC;
    AXI_11_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_11_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_11_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_11_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_11_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_11_AWVALID : IN STD_LOGIC;
    AXI_11_RREADY : IN STD_LOGIC;
    AXI_11_BREADY : IN STD_LOGIC;
    AXI_11_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_11_WLAST : IN STD_LOGIC;
    AXI_11_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_11_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_11_WVALID : IN STD_LOGIC;
    AXI_12_ACLK : IN STD_LOGIC;
    AXI_12_ARESET_N : IN STD_LOGIC;
    AXI_12_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_12_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_12_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_12_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_12_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_12_ARVALID : IN STD_LOGIC;
    AXI_12_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_12_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_12_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_12_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_12_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_12_AWVALID : IN STD_LOGIC;
    AXI_12_RREADY : IN STD_LOGIC;
    AXI_12_BREADY : IN STD_LOGIC;
    AXI_12_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_12_WLAST : IN STD_LOGIC;
    AXI_12_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_12_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_12_WVALID : IN STD_LOGIC;
    AXI_13_ACLK : IN STD_LOGIC;
    AXI_13_ARESET_N : IN STD_LOGIC;
    AXI_13_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_13_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_13_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_13_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_13_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_13_ARVALID : IN STD_LOGIC;
    AXI_13_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_13_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_13_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_13_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_13_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_13_AWVALID : IN STD_LOGIC;
    AXI_13_RREADY : IN STD_LOGIC;
    AXI_13_BREADY : IN STD_LOGIC;
    AXI_13_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_13_WLAST : IN STD_LOGIC;
    AXI_13_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_13_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_13_WVALID : IN STD_LOGIC;
    AXI_14_ACLK : IN STD_LOGIC;
    AXI_14_ARESET_N : IN STD_LOGIC;
    AXI_14_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_14_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_14_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_14_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_14_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_14_ARVALID : IN STD_LOGIC;
    AXI_14_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_14_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_14_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_14_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_14_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_14_AWVALID : IN STD_LOGIC;
    AXI_14_RREADY : IN STD_LOGIC;
    AXI_14_BREADY : IN STD_LOGIC;
    AXI_14_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_14_WLAST : IN STD_LOGIC;
    AXI_14_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_14_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_14_WVALID : IN STD_LOGIC;
    AXI_15_ACLK : IN STD_LOGIC;
    AXI_15_ARESET_N : IN STD_LOGIC;
    AXI_15_ARADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_15_ARBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_15_ARID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_15_ARLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_15_ARSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_15_ARVALID : IN STD_LOGIC;
    AXI_15_AWADDR : IN STD_LOGIC_VECTOR(32 DOWNTO 0);
    AXI_15_AWBURST : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_15_AWID : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_15_AWLEN : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    AXI_15_AWSIZE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    AXI_15_AWVALID : IN STD_LOGIC;
    AXI_15_RREADY : IN STD_LOGIC;
    AXI_15_BREADY : IN STD_LOGIC;
    AXI_15_WDATA : IN STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_15_WLAST : IN STD_LOGIC;
    AXI_15_WSTRB : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_15_WDATA_PARITY : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_15_WVALID : IN STD_LOGIC;
    APB_0_PWDATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    APB_0_PADDR : IN STD_LOGIC_VECTOR(21 DOWNTO 0);
    APB_0_PCLK : IN STD_LOGIC;
    APB_0_PENABLE : IN STD_LOGIC;
    APB_0_PRESET_N : IN STD_LOGIC;
    APB_0_PSEL : IN STD_LOGIC;
    APB_0_PWRITE : IN STD_LOGIC;
    AXI_00_ARREADY : OUT STD_LOGIC;
    AXI_00_AWREADY : OUT STD_LOGIC;
    AXI_00_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_00_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_00_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_00_RLAST : OUT STD_LOGIC;
    AXI_00_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_00_RVALID : OUT STD_LOGIC;
    AXI_00_WREADY : OUT STD_LOGIC;
    AXI_00_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_00_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_00_BVALID : OUT STD_LOGIC;
    AXI_01_ARREADY : OUT STD_LOGIC;
    AXI_01_AWREADY : OUT STD_LOGIC;
    AXI_01_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_01_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_01_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_01_RLAST : OUT STD_LOGIC;
    AXI_01_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_01_RVALID : OUT STD_LOGIC;
    AXI_01_WREADY : OUT STD_LOGIC;
    AXI_01_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_01_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_01_BVALID : OUT STD_LOGIC;
    AXI_02_ARREADY : OUT STD_LOGIC;
    AXI_02_AWREADY : OUT STD_LOGIC;
    AXI_02_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_02_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_02_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_02_RLAST : OUT STD_LOGIC;
    AXI_02_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_02_RVALID : OUT STD_LOGIC;
    AXI_02_WREADY : OUT STD_LOGIC;
    AXI_02_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_02_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_02_BVALID : OUT STD_LOGIC;
    AXI_03_ARREADY : OUT STD_LOGIC;
    AXI_03_AWREADY : OUT STD_LOGIC;
    AXI_03_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_03_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_03_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_03_RLAST : OUT STD_LOGIC;
    AXI_03_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_03_RVALID : OUT STD_LOGIC;
    AXI_03_WREADY : OUT STD_LOGIC;
    AXI_03_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_03_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_03_BVALID : OUT STD_LOGIC;
    AXI_04_ARREADY : OUT STD_LOGIC;
    AXI_04_AWREADY : OUT STD_LOGIC;
    AXI_04_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_04_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_04_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_04_RLAST : OUT STD_LOGIC;
    AXI_04_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_04_RVALID : OUT STD_LOGIC;
    AXI_04_WREADY : OUT STD_LOGIC;
    AXI_04_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_04_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_04_BVALID : OUT STD_LOGIC;
    AXI_05_ARREADY : OUT STD_LOGIC;
    AXI_05_AWREADY : OUT STD_LOGIC;
    AXI_05_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_05_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_05_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_05_RLAST : OUT STD_LOGIC;
    AXI_05_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_05_RVALID : OUT STD_LOGIC;
    AXI_05_WREADY : OUT STD_LOGIC;
    AXI_05_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_05_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_05_BVALID : OUT STD_LOGIC;
    AXI_06_ARREADY : OUT STD_LOGIC;
    AXI_06_AWREADY : OUT STD_LOGIC;
    AXI_06_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_06_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_06_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_06_RLAST : OUT STD_LOGIC;
    AXI_06_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_06_RVALID : OUT STD_LOGIC;
    AXI_06_WREADY : OUT STD_LOGIC;
    AXI_06_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_06_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_06_BVALID : OUT STD_LOGIC;
    AXI_07_ARREADY : OUT STD_LOGIC;
    AXI_07_AWREADY : OUT STD_LOGIC;
    AXI_07_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_07_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_07_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_07_RLAST : OUT STD_LOGIC;
    AXI_07_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_07_RVALID : OUT STD_LOGIC;
    AXI_07_WREADY : OUT STD_LOGIC;
    AXI_07_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_07_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_07_BVALID : OUT STD_LOGIC;
    AXI_08_ARREADY : OUT STD_LOGIC;
    AXI_08_AWREADY : OUT STD_LOGIC;
    AXI_08_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_08_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_08_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_08_RLAST : OUT STD_LOGIC;
    AXI_08_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_08_RVALID : OUT STD_LOGIC;
    AXI_08_WREADY : OUT STD_LOGIC;
    AXI_08_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_08_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_08_BVALID : OUT STD_LOGIC;
    AXI_09_ARREADY : OUT STD_LOGIC;
    AXI_09_AWREADY : OUT STD_LOGIC;
    AXI_09_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_09_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_09_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_09_RLAST : OUT STD_LOGIC;
    AXI_09_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_09_RVALID : OUT STD_LOGIC;
    AXI_09_WREADY : OUT STD_LOGIC;
    AXI_09_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_09_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_09_BVALID : OUT STD_LOGIC;
    AXI_10_ARREADY : OUT STD_LOGIC;
    AXI_10_AWREADY : OUT STD_LOGIC;
    AXI_10_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_10_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_10_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_10_RLAST : OUT STD_LOGIC;
    AXI_10_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_10_RVALID : OUT STD_LOGIC;
    AXI_10_WREADY : OUT STD_LOGIC;
    AXI_10_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_10_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_10_BVALID : OUT STD_LOGIC;
    AXI_11_ARREADY : OUT STD_LOGIC;
    AXI_11_AWREADY : OUT STD_LOGIC;
    AXI_11_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_11_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_11_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_11_RLAST : OUT STD_LOGIC;
    AXI_11_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_11_RVALID : OUT STD_LOGIC;
    AXI_11_WREADY : OUT STD_LOGIC;
    AXI_11_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_11_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_11_BVALID : OUT STD_LOGIC;
    AXI_12_ARREADY : OUT STD_LOGIC;
    AXI_12_AWREADY : OUT STD_LOGIC;
    AXI_12_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_12_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_12_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_12_RLAST : OUT STD_LOGIC;
    AXI_12_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_12_RVALID : OUT STD_LOGIC;
    AXI_12_WREADY : OUT STD_LOGIC;
    AXI_12_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_12_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_12_BVALID : OUT STD_LOGIC;
    AXI_13_ARREADY : OUT STD_LOGIC;
    AXI_13_AWREADY : OUT STD_LOGIC;
    AXI_13_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_13_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_13_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_13_RLAST : OUT STD_LOGIC;
    AXI_13_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_13_RVALID : OUT STD_LOGIC;
    AXI_13_WREADY : OUT STD_LOGIC;
    AXI_13_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_13_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_13_BVALID : OUT STD_LOGIC;
    AXI_14_ARREADY : OUT STD_LOGIC;
    AXI_14_AWREADY : OUT STD_LOGIC;
    AXI_14_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_14_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_14_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_14_RLAST : OUT STD_LOGIC;
    AXI_14_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_14_RVALID : OUT STD_LOGIC;
    AXI_14_WREADY : OUT STD_LOGIC;
    AXI_14_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_14_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_14_BVALID : OUT STD_LOGIC;
    AXI_15_ARREADY : OUT STD_LOGIC;
    AXI_15_AWREADY : OUT STD_LOGIC;
    AXI_15_RDATA_PARITY : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    AXI_15_RDATA : OUT STD_LOGIC_VECTOR(255 DOWNTO 0);
    AXI_15_RID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_15_RLAST : OUT STD_LOGIC;
    AXI_15_RRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_15_RVALID : OUT STD_LOGIC;
    AXI_15_WREADY : OUT STD_LOGIC;
    AXI_15_BID : OUT STD_LOGIC_VECTOR(5 DOWNTO 0);
    AXI_15_BRESP : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    AXI_15_BVALID : OUT STD_LOGIC;
    APB_0_PRDATA : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    APB_0_PREADY : OUT STD_LOGIC;
    APB_0_PSLVERR : OUT STD_LOGIC;
    apb_complete_0 : OUT STD_LOGIC;
    DRAM_0_STAT_CATTRIP : OUT STD_LOGIC;
    DRAM_0_STAT_TEMP : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
  );
END COMPONENT;



END tech_hbm_component_pkg;

