-------------------------------------------------------------------------------
--
-- File Name: kcu105_board_pkg.vhd
-- Contributing Authors: Andrew Brown
-- Type: RTL
-- Created: Tuesday Nov 28 16:40:00 2017
-- Template Rev: 1.0
--
-- Title: KCU105 Board Library Defines
--
-- Description:
--
--
-- Compiler options:
--
--
-- Dependencies:
--
--
--
-------------------------------------------------------------------------------

LIBRARY IEEE, common_lib;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE common_lib.common_pkg.ALL;

PACKAGE board_pkg IS



END board_pkg;
