LIBRARY IEEE, technology_lib;
USE IEEE.std_logic_1164.ALL;
USE technology_lib.technology_pkg.ALL;


PACKAGE tech_mac_10g_quad_pkg IS

   TYPE t_quad_locations_10g IS (
      QUAD_10G_122, QUAD_10G_124, QUAD_10G_125, QUAD_10G_126, QUAD_10G_131, QUAD_10G_130, QUAD_10G_128);


END tech_mac_10g_quad_pkg;

