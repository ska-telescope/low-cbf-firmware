
-------------------------------------------------------------------------------
-- (c) Copyright - Commonwealth Scientific and Industrial Research Organisation
-- (CSIRO) - 2017
--
-- All Rights Reserved.
--
-- Restricted Use.
--
-- Copyright protects this code. Except as permitted by the Copyright Act, you
-- may only use the code as expressly permitted under the terms on which the
-- code was licensed to you.
--
-------------------------------------------------------------------------------
--
-- File Name: CSIRO_ASKAP_VHDL_template.vhd
-- Contributing Authors:
-- Type: RTL
-- Created: Wed Jul 29 09:28:08 2009
-- Template Rev: 1.0
--
-- Title: (Short Description) Template file for VHDL source code for the SKA Low CBF
-- project.
--
-- Description:
--
--
--
-- Compiler options:
-- 
-- 
-- Dependencies:
-- 
-- 
-- 
-------------------------------------------------------------------------------

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;



-------------------------------------------------------------------------------
ENTITY <entity_name> IS
  PORT (

    );
END <entity_name>;

-------------------------------------------------------------------------------
ARCHITECTURE rtl OF <entity_name> IS


  ---------------------------------------------------------------------------
  -- CONSTANT, TYPE AND GENERIC DEFINITIONS  --
  ---------------------------------------------------------------------------


  ---------------------------------------------------------------------------
  -- SIGNAL DECLARATIONS  --
  ---------------------------------------------------------------------------


  ---------------------------------------------------------------------------
  -- COMPONENT DECLARATIONS  --
  ---------------------------------------------------------------------------



BEGIN


  ---------------------------------------------------------------------------
  -- INSTANTIATE COMPONENTS  --
  ---------------------------------------------------------------------------


  ---------------------------------------------------------------------------
  -- CONCURRENT SIGNAL ASSIGNMENTS  --
  ---------------------------------------------------------------------------


  ---------------------------------------------------------------------------
  -- CONCURRENT PROCESSES  --
  ---------------------------------------------------------------------------

  ---------------------------------------------------------------------------
  -- Process: <entity_name>_PROCESS
  -- Purpose:
  -- Inputs:
  -- Outputs:
  ---------------------------------------------------------------------------
  <entity_name>_process : PROCESS
                 
  BEGIN

  END PROCESS;  --  <entity_name>_process;

END rtl;
-------------------------------------------------------------------------------



