LIBRARY IEEE, technology_lib, common_lib;
USE IEEE.std_logic_1164.ALL;
USE common_lib.common_pkg.ALL;
USE common_lib.common_interface_layers_pkg.ALL;
USE technology_lib.technology_pkg.ALL;


PACKAGE tech_mac_10g_quad_component_pkg IS

COMPONENT mac_10g_quad_122
  PORT (
    gt_rxp_in_0 : IN STD_LOGIC;
    gt_rxp_in_1 : IN STD_LOGIC;
    gt_rxp_in_2 : IN STD_LOGIC;
    gt_rxp_in_3 : IN STD_LOGIC;
    gt_rxn_in_0 : IN STD_LOGIC;
    gt_rxn_in_1 : IN STD_LOGIC;
    gt_rxn_in_2 : IN STD_LOGIC;
    gt_rxn_in_3 : IN STD_LOGIC;
    gt_txp_out_0 : OUT STD_LOGIC;
    gt_txp_out_1 : OUT STD_LOGIC;
    gt_txp_out_2 : OUT STD_LOGIC;
    gt_txp_out_3 : OUT STD_LOGIC;
    gt_txn_out_0 : OUT STD_LOGIC;
    gt_txn_out_1 : OUT STD_LOGIC;
    gt_txn_out_2 : OUT STD_LOGIC;
    gt_txn_out_3 : OUT STD_LOGIC;
    rx_core_clk_0 : IN STD_LOGIC;
    rx_core_clk_1 : IN STD_LOGIC;
    rx_core_clk_2 : IN STD_LOGIC;
    rx_core_clk_3 : IN STD_LOGIC;
    txoutclksel_in_0 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    rxoutclksel_in_0 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    txoutclksel_in_1 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    rxoutclksel_in_1 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    txoutclksel_in_2 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    rxoutclksel_in_2 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    txoutclksel_in_3 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    rxoutclksel_in_3 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    gt_dmonitorout_0 : OUT STD_LOGIC_VECTOR(16 DOWNTO 0);
    gt_dmonitorout_1 : OUT STD_LOGIC_VECTOR(16 DOWNTO 0);
    gt_dmonitorout_2 : OUT STD_LOGIC_VECTOR(16 DOWNTO 0);
    gt_dmonitorout_3 : OUT STD_LOGIC_VECTOR(16 DOWNTO 0);
    gt_eyescandataerror_0 : OUT STD_LOGIC;
    gt_eyescandataerror_1 : OUT STD_LOGIC;
    gt_eyescandataerror_2 : OUT STD_LOGIC;
    gt_eyescandataerror_3 : OUT STD_LOGIC;
    gt_eyescanreset_0 : IN STD_LOGIC;
    gt_eyescanreset_1 : IN STD_LOGIC;
    gt_eyescanreset_2 : IN STD_LOGIC;
    gt_eyescanreset_3 : IN STD_LOGIC;
    gt_eyescantrigger_0 : IN STD_LOGIC;
    gt_eyescantrigger_1 : IN STD_LOGIC;
    gt_eyescantrigger_2 : IN STD_LOGIC;
    gt_eyescantrigger_3 : IN STD_LOGIC;
    gt_pcsrsvdin_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_pcsrsvdin_1 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_pcsrsvdin_2 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_pcsrsvdin_3 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_rxbufreset_0 : IN STD_LOGIC;
    gt_rxbufreset_1 : IN STD_LOGIC;
    gt_rxbufreset_2 : IN STD_LOGIC;
    gt_rxbufreset_3 : IN STD_LOGIC;
    gt_rxbufstatus_0 : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
    gt_rxbufstatus_1 : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
    gt_rxbufstatus_2 : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
    gt_rxbufstatus_3 : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
    gt_rxcdrhold_0 : IN STD_LOGIC;
    gt_rxcdrhold_1 : IN STD_LOGIC;
    gt_rxcdrhold_2 : IN STD_LOGIC;
    gt_rxcdrhold_3 : IN STD_LOGIC;
    gt_rxcommadeten_0 : IN STD_LOGIC;
    gt_rxcommadeten_1 : IN STD_LOGIC;
    gt_rxcommadeten_2 : IN STD_LOGIC;
    gt_rxcommadeten_3 : IN STD_LOGIC;
    gt_rxdfeagchold_0 : IN STD_LOGIC;
    gt_rxdfeagchold_1 : IN STD_LOGIC;
    gt_rxdfeagchold_2 : IN STD_LOGIC;
    gt_rxdfeagchold_3 : IN STD_LOGIC;
    gt_rxdfelpmreset_0 : IN STD_LOGIC;
    gt_rxdfelpmreset_1 : IN STD_LOGIC;
    gt_rxdfelpmreset_2 : IN STD_LOGIC;
    gt_rxdfelpmreset_3 : IN STD_LOGIC;
    gt_rxlatclk_0 : IN STD_LOGIC;
    gt_rxlatclk_1 : IN STD_LOGIC;
    gt_rxlatclk_2 : IN STD_LOGIC;
    gt_rxlatclk_3 : IN STD_LOGIC;
    gt_rxlpmen_0 : IN STD_LOGIC;
    gt_rxlpmen_1 : IN STD_LOGIC;
    gt_rxlpmen_2 : IN STD_LOGIC;
    gt_rxlpmen_3 : IN STD_LOGIC;
    gt_rxpcsreset_0 : IN STD_LOGIC;
    gt_rxpcsreset_1 : IN STD_LOGIC;
    gt_rxpcsreset_2 : IN STD_LOGIC;
    gt_rxpcsreset_3 : IN STD_LOGIC;
    gt_rxpmareset_0 : IN STD_LOGIC;
    gt_rxpmareset_1 : IN STD_LOGIC;
    gt_rxpmareset_2 : IN STD_LOGIC;
    gt_rxpmareset_3 : IN STD_LOGIC;
    gt_rxpolarity_0 : IN STD_LOGIC;
    gt_rxpolarity_1 : IN STD_LOGIC;
    gt_rxpolarity_2 : IN STD_LOGIC;
    gt_rxpolarity_3 : IN STD_LOGIC;
    gt_rxprbscntreset_0 : IN STD_LOGIC;
    gt_rxprbscntreset_1 : IN STD_LOGIC;
    gt_rxprbscntreset_2 : IN STD_LOGIC;
    gt_rxprbscntreset_3 : IN STD_LOGIC;
    gt_rxprbserr_0 : OUT STD_LOGIC;
    gt_rxprbserr_1 : OUT STD_LOGIC;
    gt_rxprbserr_2 : OUT STD_LOGIC;
    gt_rxprbserr_3 : OUT STD_LOGIC;
    gt_rxprbssel_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbssel_1 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbssel_2 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxprbssel_3 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_rxrate_0 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    gt_rxrate_1 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    gt_rxrate_2 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    gt_rxrate_3 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    gt_rxslide_in_0 : IN STD_LOGIC;
    gt_rxslide_in_1 : IN STD_LOGIC;
    gt_rxslide_in_2 : IN STD_LOGIC;
    gt_rxslide_in_3 : IN STD_LOGIC;
    gt_rxstartofseq_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    gt_rxstartofseq_1 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    gt_rxstartofseq_2 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    gt_rxstartofseq_3 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    gt_txbufstatus_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    gt_txbufstatus_1 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    gt_txbufstatus_2 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    gt_txbufstatus_3 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    gt_txdiffctrl_0 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    gt_txdiffctrl_1 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    gt_txdiffctrl_2 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    gt_txdiffctrl_3 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    gt_txinhibit_0 : IN STD_LOGIC;
    gt_txinhibit_1 : IN STD_LOGIC;
    gt_txinhibit_2 : IN STD_LOGIC;
    gt_txinhibit_3 : IN STD_LOGIC;
    gt_txlatclk_0 : IN STD_LOGIC;
    gt_txlatclk_1 : IN STD_LOGIC;
    gt_txlatclk_2 : IN STD_LOGIC;
    gt_txlatclk_3 : IN STD_LOGIC;
    gt_txmaincursor_0 : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    gt_txmaincursor_1 : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    gt_txmaincursor_2 : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    gt_txmaincursor_3 : IN STD_LOGIC_VECTOR(6 DOWNTO 0);
    gt_txpcsreset_0 : IN STD_LOGIC;
    gt_txpcsreset_1 : IN STD_LOGIC;
    gt_txpcsreset_2 : IN STD_LOGIC;
    gt_txpcsreset_3 : IN STD_LOGIC;
    gt_txpmareset_0 : IN STD_LOGIC;
    gt_txpmareset_1 : IN STD_LOGIC;
    gt_txpmareset_2 : IN STD_LOGIC;
    gt_txpmareset_3 : IN STD_LOGIC;
    gt_txpolarity_0 : IN STD_LOGIC;
    gt_txpolarity_1 : IN STD_LOGIC;
    gt_txpolarity_2 : IN STD_LOGIC;
    gt_txpolarity_3 : IN STD_LOGIC;
    gt_txpostcursor_0 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    gt_txpostcursor_1 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    gt_txpostcursor_2 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    gt_txpostcursor_3 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    gt_txprbsforceerr_0 : IN STD_LOGIC;
    gt_txprbsforceerr_1 : IN STD_LOGIC;
    gt_txprbsforceerr_2 : IN STD_LOGIC;
    gt_txprbsforceerr_3 : IN STD_LOGIC;
    gt_txprbssel_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txprbssel_1 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txprbssel_2 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txprbssel_3 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    gt_txprecursor_0 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    gt_txprecursor_1 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    gt_txprecursor_2 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    gt_txprecursor_3 : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
    gtwiz_reset_tx_datapath_0 : IN STD_LOGIC;
    gtwiz_reset_tx_datapath_1 : IN STD_LOGIC;
    gtwiz_reset_tx_datapath_2 : IN STD_LOGIC;
    gtwiz_reset_tx_datapath_3 : IN STD_LOGIC;
    gtwiz_reset_rx_datapath_0 : IN STD_LOGIC;
    gtwiz_reset_rx_datapath_1 : IN STD_LOGIC;
    gtwiz_reset_rx_datapath_2 : IN STD_LOGIC;
    gtwiz_reset_rx_datapath_3 : IN STD_LOGIC;
    rxrecclkout_0 : OUT STD_LOGIC;
    rxrecclkout_1 : OUT STD_LOGIC;
    rxrecclkout_2 : OUT STD_LOGIC;
    rxrecclkout_3 : OUT STD_LOGIC;
    gt_drpclk_0 : IN STD_LOGIC;
    gt_drpclk_1 : IN STD_LOGIC;
    gt_drpclk_2 : IN STD_LOGIC;
    gt_drpclk_3 : IN STD_LOGIC;
    gt_drpdo_0 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_drpdo_1 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_drpdo_2 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_drpdo_3 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_drprdy_0 : OUT STD_LOGIC;
    gt_drprdy_1 : OUT STD_LOGIC;
    gt_drprdy_2 : OUT STD_LOGIC;
    gt_drprdy_3 : OUT STD_LOGIC;
    gt_drpen_0 : IN STD_LOGIC;
    gt_drpen_1 : IN STD_LOGIC;
    gt_drpen_2 : IN STD_LOGIC;
    gt_drpen_3 : IN STD_LOGIC;
    gt_drpwe_0 : IN STD_LOGIC;
    gt_drpwe_1 : IN STD_LOGIC;
    gt_drpwe_2 : IN STD_LOGIC;
    gt_drpwe_3 : IN STD_LOGIC;
    gt_drpaddr_0 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_drpaddr_1 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_drpaddr_2 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_drpaddr_3 : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
    gt_drpdi_0 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_drpdi_1 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_drpdi_2 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    gt_drpdi_3 : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
    sys_reset : IN STD_LOGIC;
    dclk : IN STD_LOGIC;
    tx_clk_out_0 : OUT STD_LOGIC;
    tx_clk_out_1 : OUT STD_LOGIC;
    tx_clk_out_2 : OUT STD_LOGIC;
    tx_clk_out_3 : OUT STD_LOGIC;
    rx_clk_out_0 : OUT STD_LOGIC;
    rx_clk_out_1 : OUT STD_LOGIC;
    rx_clk_out_2 : OUT STD_LOGIC;
    rx_clk_out_3 : OUT STD_LOGIC;
    gt_refclk_p : IN STD_LOGIC;
    gt_refclk_n : IN STD_LOGIC;
    gt_refclk_out : OUT STD_LOGIC;
    gtpowergood_out_0 : OUT STD_LOGIC;
    gtpowergood_out_1 : OUT STD_LOGIC;
    gtpowergood_out_2 : OUT STD_LOGIC;
    gtpowergood_out_3 : OUT STD_LOGIC;
    rx_reset_0 : IN STD_LOGIC;
    rx_reset_1 : IN STD_LOGIC;
    rx_reset_2 : IN STD_LOGIC;
    rx_reset_3 : IN STD_LOGIC;
    user_rx_reset_0 : OUT STD_LOGIC;
    user_rx_reset_1 : OUT STD_LOGIC;
    user_rx_reset_2 : OUT STD_LOGIC;
    user_rx_reset_3 : OUT STD_LOGIC;
    rx_axis_tvalid_0 : OUT STD_LOGIC;
    rx_axis_tvalid_1 : OUT STD_LOGIC;
    rx_axis_tvalid_2 : OUT STD_LOGIC;
    rx_axis_tvalid_3 : OUT STD_LOGIC;
    rx_axis_tdata_0 : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
    rx_axis_tdata_1 : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
    rx_axis_tdata_2 : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
    rx_axis_tdata_3 : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
    rx_axis_tlast_0 : OUT STD_LOGIC;
    rx_axis_tlast_1 : OUT STD_LOGIC;
    rx_axis_tlast_2 : OUT STD_LOGIC;
    rx_axis_tlast_3 : OUT STD_LOGIC;
    rx_axis_tkeep_0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    rx_axis_tkeep_1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    rx_axis_tkeep_2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    rx_axis_tkeep_3 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    rx_axis_tuser_0 : OUT STD_LOGIC;
    rx_axis_tuser_1 : OUT STD_LOGIC;
    rx_axis_tuser_2 : OUT STD_LOGIC;
    rx_axis_tuser_3 : OUT STD_LOGIC;
    ctl_rx_enable_0 : IN STD_LOGIC;
    ctl_rx_enable_1 : IN STD_LOGIC;
    ctl_rx_enable_2 : IN STD_LOGIC;
    ctl_rx_enable_3 : IN STD_LOGIC;
    ctl_rx_check_preamble_0 : IN STD_LOGIC;
    ctl_rx_check_preamble_1 : IN STD_LOGIC;
    ctl_rx_check_preamble_2 : IN STD_LOGIC;
    ctl_rx_check_preamble_3 : IN STD_LOGIC;
    ctl_rx_check_sfd_0 : IN STD_LOGIC;
    ctl_rx_check_sfd_1 : IN STD_LOGIC;
    ctl_rx_check_sfd_2 : IN STD_LOGIC;
    ctl_rx_check_sfd_3 : IN STD_LOGIC;
    ctl_rx_force_resync_0 : IN STD_LOGIC;
    ctl_rx_force_resync_1 : IN STD_LOGIC;
    ctl_rx_force_resync_2 : IN STD_LOGIC;
    ctl_rx_force_resync_3 : IN STD_LOGIC;
    ctl_rx_delete_fcs_0 : IN STD_LOGIC;
    ctl_rx_delete_fcs_1 : IN STD_LOGIC;
    ctl_rx_delete_fcs_2 : IN STD_LOGIC;
    ctl_rx_delete_fcs_3 : IN STD_LOGIC;
    ctl_rx_ignore_fcs_0 : IN STD_LOGIC;
    ctl_rx_ignore_fcs_1 : IN STD_LOGIC;
    ctl_rx_ignore_fcs_2 : IN STD_LOGIC;
    ctl_rx_ignore_fcs_3 : IN STD_LOGIC;
    ctl_rx_max_packet_len_0 : IN STD_LOGIC_VECTOR(14 DOWNTO 0);
    ctl_rx_max_packet_len_1 : IN STD_LOGIC_VECTOR(14 DOWNTO 0);
    ctl_rx_max_packet_len_2 : IN STD_LOGIC_VECTOR(14 DOWNTO 0);
    ctl_rx_max_packet_len_3 : IN STD_LOGIC_VECTOR(14 DOWNTO 0);
    ctl_rx_min_packet_len_0 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    ctl_rx_min_packet_len_1 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    ctl_rx_min_packet_len_2 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    ctl_rx_min_packet_len_3 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    ctl_rx_process_lfi_0 : IN STD_LOGIC;
    ctl_rx_process_lfi_1 : IN STD_LOGIC;
    ctl_rx_process_lfi_2 : IN STD_LOGIC;
    ctl_rx_process_lfi_3 : IN STD_LOGIC;
    ctl_rx_test_pattern_0 : IN STD_LOGIC;
    ctl_rx_test_pattern_1 : IN STD_LOGIC;
    ctl_rx_test_pattern_2 : IN STD_LOGIC;
    ctl_rx_test_pattern_3 : IN STD_LOGIC;
    ctl_rx_data_pattern_select_0 : IN STD_LOGIC;
    ctl_rx_data_pattern_select_1 : IN STD_LOGIC;
    ctl_rx_data_pattern_select_2 : IN STD_LOGIC;
    ctl_rx_data_pattern_select_3 : IN STD_LOGIC;
    ctl_rx_test_pattern_enable_0 : IN STD_LOGIC;
    ctl_rx_test_pattern_enable_1 : IN STD_LOGIC;
    ctl_rx_test_pattern_enable_2 : IN STD_LOGIC;
    ctl_rx_test_pattern_enable_3 : IN STD_LOGIC;
    ctl_rx_custom_preamble_enable_0 : IN STD_LOGIC;
    ctl_rx_custom_preamble_enable_1 : IN STD_LOGIC;
    ctl_rx_custom_preamble_enable_2 : IN STD_LOGIC;
    ctl_rx_custom_preamble_enable_3 : IN STD_LOGIC;
    stat_rx_framing_err_0 : OUT STD_LOGIC;
    stat_rx_framing_err_1 : OUT STD_LOGIC;
    stat_rx_framing_err_2 : OUT STD_LOGIC;
    stat_rx_framing_err_3 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_0 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_1 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_2 : OUT STD_LOGIC;
    stat_rx_framing_err_valid_3 : OUT STD_LOGIC;
    stat_rx_local_fault_0 : OUT STD_LOGIC;
    stat_rx_local_fault_1 : OUT STD_LOGIC;
    stat_rx_local_fault_2 : OUT STD_LOGIC;
    stat_rx_local_fault_3 : OUT STD_LOGIC;
    stat_rx_block_lock_0 : OUT STD_LOGIC;
    stat_rx_block_lock_1 : OUT STD_LOGIC;
    stat_rx_block_lock_2 : OUT STD_LOGIC;
    stat_rx_block_lock_3 : OUT STD_LOGIC;
    stat_rx_valid_ctrl_code_0 : OUT STD_LOGIC;
    stat_rx_valid_ctrl_code_1 : OUT STD_LOGIC;
    stat_rx_valid_ctrl_code_2 : OUT STD_LOGIC;
    stat_rx_valid_ctrl_code_3 : OUT STD_LOGIC;
    stat_rx_status_0 : OUT STD_LOGIC;
    stat_rx_status_1 : OUT STD_LOGIC;
    stat_rx_status_2 : OUT STD_LOGIC;
    stat_rx_status_3 : OUT STD_LOGIC;
    stat_rx_remote_fault_0 : OUT STD_LOGIC;
    stat_rx_remote_fault_1 : OUT STD_LOGIC;
    stat_rx_remote_fault_2 : OUT STD_LOGIC;
    stat_rx_remote_fault_3 : OUT STD_LOGIC;
    stat_rx_bad_fcs_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_bad_fcs_1 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_bad_fcs_2 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_bad_fcs_3 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_stomped_fcs_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_stomped_fcs_1 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_stomped_fcs_2 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_stomped_fcs_3 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_truncated_0 : OUT STD_LOGIC;
    stat_rx_truncated_1 : OUT STD_LOGIC;
    stat_rx_truncated_2 : OUT STD_LOGIC;
    stat_rx_truncated_3 : OUT STD_LOGIC;
    stat_rx_internal_local_fault_0 : OUT STD_LOGIC;
    stat_rx_internal_local_fault_1 : OUT STD_LOGIC;
    stat_rx_internal_local_fault_2 : OUT STD_LOGIC;
    stat_rx_internal_local_fault_3 : OUT STD_LOGIC;
    stat_rx_received_local_fault_0 : OUT STD_LOGIC;
    stat_rx_received_local_fault_1 : OUT STD_LOGIC;
    stat_rx_received_local_fault_2 : OUT STD_LOGIC;
    stat_rx_received_local_fault_3 : OUT STD_LOGIC;
    stat_rx_hi_ber_0 : OUT STD_LOGIC;
    stat_rx_hi_ber_1 : OUT STD_LOGIC;
    stat_rx_hi_ber_2 : OUT STD_LOGIC;
    stat_rx_hi_ber_3 : OUT STD_LOGIC;
    stat_rx_got_signal_os_0 : OUT STD_LOGIC;
    stat_rx_got_signal_os_1 : OUT STD_LOGIC;
    stat_rx_got_signal_os_2 : OUT STD_LOGIC;
    stat_rx_got_signal_os_3 : OUT STD_LOGIC;
    stat_rx_test_pattern_mismatch_0 : OUT STD_LOGIC;
    stat_rx_test_pattern_mismatch_1 : OUT STD_LOGIC;
    stat_rx_test_pattern_mismatch_2 : OUT STD_LOGIC;
    stat_rx_test_pattern_mismatch_3 : OUT STD_LOGIC;
    stat_rx_total_bytes_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_total_bytes_1 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_total_bytes_2 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_total_bytes_3 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_rx_total_packets_0 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_total_packets_1 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_total_packets_2 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_total_packets_3 : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    stat_rx_total_good_bytes_0 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_rx_total_good_bytes_1 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_rx_total_good_bytes_2 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_rx_total_good_bytes_3 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_rx_total_good_packets_0 : OUT STD_LOGIC;
    stat_rx_total_good_packets_1 : OUT STD_LOGIC;
    stat_rx_total_good_packets_2 : OUT STD_LOGIC;
    stat_rx_total_good_packets_3 : OUT STD_LOGIC;
    stat_rx_packet_bad_fcs_0 : OUT STD_LOGIC;
    stat_rx_packet_bad_fcs_1 : OUT STD_LOGIC;
    stat_rx_packet_bad_fcs_2 : OUT STD_LOGIC;
    stat_rx_packet_bad_fcs_3 : OUT STD_LOGIC;
    stat_rx_packet_64_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_64_bytes_1 : OUT STD_LOGIC;
    stat_rx_packet_64_bytes_2 : OUT STD_LOGIC;
    stat_rx_packet_64_bytes_3 : OUT STD_LOGIC;
    stat_rx_packet_65_127_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_65_127_bytes_1 : OUT STD_LOGIC;
    stat_rx_packet_65_127_bytes_2 : OUT STD_LOGIC;
    stat_rx_packet_65_127_bytes_3 : OUT STD_LOGIC;
    stat_rx_packet_128_255_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_128_255_bytes_1 : OUT STD_LOGIC;
    stat_rx_packet_128_255_bytes_2 : OUT STD_LOGIC;
    stat_rx_packet_128_255_bytes_3 : OUT STD_LOGIC;
    stat_rx_packet_256_511_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_256_511_bytes_1 : OUT STD_LOGIC;
    stat_rx_packet_256_511_bytes_2 : OUT STD_LOGIC;
    stat_rx_packet_256_511_bytes_3 : OUT STD_LOGIC;
    stat_rx_packet_512_1023_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_512_1023_bytes_1 : OUT STD_LOGIC;
    stat_rx_packet_512_1023_bytes_2 : OUT STD_LOGIC;
    stat_rx_packet_512_1023_bytes_3 : OUT STD_LOGIC;
    stat_rx_packet_1024_1518_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1024_1518_bytes_1 : OUT STD_LOGIC;
    stat_rx_packet_1024_1518_bytes_2 : OUT STD_LOGIC;
    stat_rx_packet_1024_1518_bytes_3 : OUT STD_LOGIC;
    stat_rx_packet_1519_1522_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1519_1522_bytes_1 : OUT STD_LOGIC;
    stat_rx_packet_1519_1522_bytes_2 : OUT STD_LOGIC;
    stat_rx_packet_1519_1522_bytes_3 : OUT STD_LOGIC;
    stat_rx_packet_1523_1548_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1523_1548_bytes_1 : OUT STD_LOGIC;
    stat_rx_packet_1523_1548_bytes_2 : OUT STD_LOGIC;
    stat_rx_packet_1523_1548_bytes_3 : OUT STD_LOGIC;
    stat_rx_packet_1549_2047_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_1549_2047_bytes_1 : OUT STD_LOGIC;
    stat_rx_packet_1549_2047_bytes_2 : OUT STD_LOGIC;
    stat_rx_packet_1549_2047_bytes_3 : OUT STD_LOGIC;
    stat_rx_packet_2048_4095_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_2048_4095_bytes_1 : OUT STD_LOGIC;
    stat_rx_packet_2048_4095_bytes_2 : OUT STD_LOGIC;
    stat_rx_packet_2048_4095_bytes_3 : OUT STD_LOGIC;
    stat_rx_packet_4096_8191_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_4096_8191_bytes_1 : OUT STD_LOGIC;
    stat_rx_packet_4096_8191_bytes_2 : OUT STD_LOGIC;
    stat_rx_packet_4096_8191_bytes_3 : OUT STD_LOGIC;
    stat_rx_packet_8192_9215_bytes_0 : OUT STD_LOGIC;
    stat_rx_packet_8192_9215_bytes_1 : OUT STD_LOGIC;
    stat_rx_packet_8192_9215_bytes_2 : OUT STD_LOGIC;
    stat_rx_packet_8192_9215_bytes_3 : OUT STD_LOGIC;
    stat_rx_packet_small_0 : OUT STD_LOGIC;
    stat_rx_packet_small_1 : OUT STD_LOGIC;
    stat_rx_packet_small_2 : OUT STD_LOGIC;
    stat_rx_packet_small_3 : OUT STD_LOGIC;
    stat_rx_packet_large_0 : OUT STD_LOGIC;
    stat_rx_packet_large_1 : OUT STD_LOGIC;
    stat_rx_packet_large_2 : OUT STD_LOGIC;
    stat_rx_packet_large_3 : OUT STD_LOGIC;
    stat_rx_oversize_0 : OUT STD_LOGIC;
    stat_rx_oversize_1 : OUT STD_LOGIC;
    stat_rx_oversize_2 : OUT STD_LOGIC;
    stat_rx_oversize_3 : OUT STD_LOGIC;
    stat_rx_toolong_0 : OUT STD_LOGIC;
    stat_rx_toolong_1 : OUT STD_LOGIC;
    stat_rx_toolong_2 : OUT STD_LOGIC;
    stat_rx_toolong_3 : OUT STD_LOGIC;
    stat_rx_undersize_0 : OUT STD_LOGIC;
    stat_rx_undersize_1 : OUT STD_LOGIC;
    stat_rx_undersize_2 : OUT STD_LOGIC;
    stat_rx_undersize_3 : OUT STD_LOGIC;
    stat_rx_fragment_0 : OUT STD_LOGIC;
    stat_rx_fragment_1 : OUT STD_LOGIC;
    stat_rx_fragment_2 : OUT STD_LOGIC;
    stat_rx_fragment_3 : OUT STD_LOGIC;
    stat_rx_jabber_0 : OUT STD_LOGIC;
    stat_rx_jabber_1 : OUT STD_LOGIC;
    stat_rx_jabber_2 : OUT STD_LOGIC;
    stat_rx_jabber_3 : OUT STD_LOGIC;
    stat_rx_bad_code_0 : OUT STD_LOGIC;
    stat_rx_bad_code_1 : OUT STD_LOGIC;
    stat_rx_bad_code_2 : OUT STD_LOGIC;
    stat_rx_bad_code_3 : OUT STD_LOGIC;
    stat_rx_bad_sfd_0 : OUT STD_LOGIC;
    stat_rx_bad_sfd_1 : OUT STD_LOGIC;
    stat_rx_bad_sfd_2 : OUT STD_LOGIC;
    stat_rx_bad_sfd_3 : OUT STD_LOGIC;
    stat_rx_bad_preamble_0 : OUT STD_LOGIC;
    stat_rx_bad_preamble_1 : OUT STD_LOGIC;
    stat_rx_bad_preamble_2 : OUT STD_LOGIC;
    stat_rx_bad_preamble_3 : OUT STD_LOGIC;
    tx_reset_0 : IN STD_LOGIC;
    tx_reset_1 : IN STD_LOGIC;
    tx_reset_2 : IN STD_LOGIC;
    tx_reset_3 : IN STD_LOGIC;
    user_tx_reset_0 : OUT STD_LOGIC;
    user_tx_reset_1 : OUT STD_LOGIC;
    user_tx_reset_2 : OUT STD_LOGIC;
    user_tx_reset_3 : OUT STD_LOGIC;
    tx_axis_tready_0 : OUT STD_LOGIC;
    tx_axis_tready_1 : OUT STD_LOGIC;
    tx_axis_tready_2 : OUT STD_LOGIC;
    tx_axis_tready_3 : OUT STD_LOGIC;
    tx_axis_tvalid_0 : IN STD_LOGIC;
    tx_axis_tvalid_1 : IN STD_LOGIC;
    tx_axis_tvalid_2 : IN STD_LOGIC;
    tx_axis_tvalid_3 : IN STD_LOGIC;
    tx_axis_tdata_0 : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
    tx_axis_tdata_1 : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
    tx_axis_tdata_2 : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
    tx_axis_tdata_3 : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
    tx_axis_tlast_0 : IN STD_LOGIC;
    tx_axis_tlast_1 : IN STD_LOGIC;
    tx_axis_tlast_2 : IN STD_LOGIC;
    tx_axis_tlast_3 : IN STD_LOGIC;
    tx_axis_tkeep_0 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    tx_axis_tkeep_1 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    tx_axis_tkeep_2 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    tx_axis_tkeep_3 : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    tx_axis_tuser_0 : IN STD_LOGIC;
    tx_axis_tuser_1 : IN STD_LOGIC;
    tx_axis_tuser_2 : IN STD_LOGIC;
    tx_axis_tuser_3 : IN STD_LOGIC;
    tx_unfout_0 : OUT STD_LOGIC;
    tx_unfout_1 : OUT STD_LOGIC;
    tx_unfout_2 : OUT STD_LOGIC;
    tx_unfout_3 : OUT STD_LOGIC;
    tx_preamblein_0 : IN STD_LOGIC_VECTOR(55 DOWNTO 0);
    rx_preambleout_0 : OUT STD_LOGIC_VECTOR(55 DOWNTO 0);
    tx_preamblein_1 : IN STD_LOGIC_VECTOR(55 DOWNTO 0);
    rx_preambleout_1 : OUT STD_LOGIC_VECTOR(55 DOWNTO 0);
    tx_preamblein_2 : IN STD_LOGIC_VECTOR(55 DOWNTO 0);
    rx_preambleout_2 : OUT STD_LOGIC_VECTOR(55 DOWNTO 0);
    tx_preamblein_3 : IN STD_LOGIC_VECTOR(55 DOWNTO 0);
    rx_preambleout_3 : OUT STD_LOGIC_VECTOR(55 DOWNTO 0);
    stat_tx_local_fault_0 : OUT STD_LOGIC;
    stat_tx_local_fault_1 : OUT STD_LOGIC;
    stat_tx_local_fault_2 : OUT STD_LOGIC;
    stat_tx_local_fault_3 : OUT STD_LOGIC;
    stat_tx_total_bytes_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_tx_total_bytes_1 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_tx_total_bytes_2 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_tx_total_bytes_3 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    stat_tx_total_packets_0 : OUT STD_LOGIC;
    stat_tx_total_packets_1 : OUT STD_LOGIC;
    stat_tx_total_packets_2 : OUT STD_LOGIC;
    stat_tx_total_packets_3 : OUT STD_LOGIC;
    stat_tx_total_good_bytes_0 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_tx_total_good_bytes_1 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_tx_total_good_bytes_2 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_tx_total_good_bytes_3 : OUT STD_LOGIC_VECTOR(13 DOWNTO 0);
    stat_tx_total_good_packets_0 : OUT STD_LOGIC;
    stat_tx_total_good_packets_1 : OUT STD_LOGIC;
    stat_tx_total_good_packets_2 : OUT STD_LOGIC;
    stat_tx_total_good_packets_3 : OUT STD_LOGIC;
    stat_tx_bad_fcs_0 : OUT STD_LOGIC;
    stat_tx_bad_fcs_1 : OUT STD_LOGIC;
    stat_tx_bad_fcs_2 : OUT STD_LOGIC;
    stat_tx_bad_fcs_3 : OUT STD_LOGIC;
    stat_tx_packet_64_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_64_bytes_1 : OUT STD_LOGIC;
    stat_tx_packet_64_bytes_2 : OUT STD_LOGIC;
    stat_tx_packet_64_bytes_3 : OUT STD_LOGIC;
    stat_tx_packet_65_127_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_65_127_bytes_1 : OUT STD_LOGIC;
    stat_tx_packet_65_127_bytes_2 : OUT STD_LOGIC;
    stat_tx_packet_65_127_bytes_3 : OUT STD_LOGIC;
    stat_tx_packet_128_255_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_128_255_bytes_1 : OUT STD_LOGIC;
    stat_tx_packet_128_255_bytes_2 : OUT STD_LOGIC;
    stat_tx_packet_128_255_bytes_3 : OUT STD_LOGIC;
    stat_tx_packet_256_511_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_256_511_bytes_1 : OUT STD_LOGIC;
    stat_tx_packet_256_511_bytes_2 : OUT STD_LOGIC;
    stat_tx_packet_256_511_bytes_3 : OUT STD_LOGIC;
    stat_tx_packet_512_1023_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_512_1023_bytes_1 : OUT STD_LOGIC;
    stat_tx_packet_512_1023_bytes_2 : OUT STD_LOGIC;
    stat_tx_packet_512_1023_bytes_3 : OUT STD_LOGIC;
    stat_tx_packet_1024_1518_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1024_1518_bytes_1 : OUT STD_LOGIC;
    stat_tx_packet_1024_1518_bytes_2 : OUT STD_LOGIC;
    stat_tx_packet_1024_1518_bytes_3 : OUT STD_LOGIC;
    stat_tx_packet_1519_1522_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1519_1522_bytes_1 : OUT STD_LOGIC;
    stat_tx_packet_1519_1522_bytes_2 : OUT STD_LOGIC;
    stat_tx_packet_1519_1522_bytes_3 : OUT STD_LOGIC;
    stat_tx_packet_1523_1548_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1523_1548_bytes_1 : OUT STD_LOGIC;
    stat_tx_packet_1523_1548_bytes_2 : OUT STD_LOGIC;
    stat_tx_packet_1523_1548_bytes_3 : OUT STD_LOGIC;
    stat_tx_packet_1549_2047_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_1549_2047_bytes_1 : OUT STD_LOGIC;
    stat_tx_packet_1549_2047_bytes_2 : OUT STD_LOGIC;
    stat_tx_packet_1549_2047_bytes_3 : OUT STD_LOGIC;
    stat_tx_packet_2048_4095_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_2048_4095_bytes_1 : OUT STD_LOGIC;
    stat_tx_packet_2048_4095_bytes_2 : OUT STD_LOGIC;
    stat_tx_packet_2048_4095_bytes_3 : OUT STD_LOGIC;
    stat_tx_packet_4096_8191_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_4096_8191_bytes_1 : OUT STD_LOGIC;
    stat_tx_packet_4096_8191_bytes_2 : OUT STD_LOGIC;
    stat_tx_packet_4096_8191_bytes_3 : OUT STD_LOGIC;
    stat_tx_packet_8192_9215_bytes_0 : OUT STD_LOGIC;
    stat_tx_packet_8192_9215_bytes_1 : OUT STD_LOGIC;
    stat_tx_packet_8192_9215_bytes_2 : OUT STD_LOGIC;
    stat_tx_packet_8192_9215_bytes_3 : OUT STD_LOGIC;
    stat_tx_packet_small_0 : OUT STD_LOGIC;
    stat_tx_packet_small_1 : OUT STD_LOGIC;
    stat_tx_packet_small_2 : OUT STD_LOGIC;
    stat_tx_packet_small_3 : OUT STD_LOGIC;
    stat_tx_packet_large_0 : OUT STD_LOGIC;
    stat_tx_packet_large_1 : OUT STD_LOGIC;
    stat_tx_packet_large_2 : OUT STD_LOGIC;
    stat_tx_packet_large_3 : OUT STD_LOGIC;
    stat_tx_frame_error_0 : OUT STD_LOGIC;
    stat_tx_frame_error_1 : OUT STD_LOGIC;
    stat_tx_frame_error_2 : OUT STD_LOGIC;
    stat_tx_frame_error_3 : OUT STD_LOGIC;
    ctl_tx_enable_0 : IN STD_LOGIC;
    ctl_tx_enable_1 : IN STD_LOGIC;
    ctl_tx_enable_2 : IN STD_LOGIC;
    ctl_tx_enable_3 : IN STD_LOGIC;
    ctl_tx_send_rfi_0 : IN STD_LOGIC;
    ctl_tx_send_rfi_1 : IN STD_LOGIC;
    ctl_tx_send_rfi_2 : IN STD_LOGIC;
    ctl_tx_send_rfi_3 : IN STD_LOGIC;
    ctl_tx_send_lfi_0 : IN STD_LOGIC;
    ctl_tx_send_lfi_1 : IN STD_LOGIC;
    ctl_tx_send_lfi_2 : IN STD_LOGIC;
    ctl_tx_send_lfi_3 : IN STD_LOGIC;
    ctl_tx_send_idle_0 : IN STD_LOGIC;
    ctl_tx_send_idle_1 : IN STD_LOGIC;
    ctl_tx_send_idle_2 : IN STD_LOGIC;
    ctl_tx_send_idle_3 : IN STD_LOGIC;
    ctl_tx_fcs_ins_enable_0 : IN STD_LOGIC;
    ctl_tx_fcs_ins_enable_1 : IN STD_LOGIC;
    ctl_tx_fcs_ins_enable_2 : IN STD_LOGIC;
    ctl_tx_fcs_ins_enable_3 : IN STD_LOGIC;
    ctl_tx_ignore_fcs_0 : IN STD_LOGIC;
    ctl_tx_ignore_fcs_1 : IN STD_LOGIC;
    ctl_tx_ignore_fcs_2 : IN STD_LOGIC;
    ctl_tx_ignore_fcs_3 : IN STD_LOGIC;
    ctl_tx_test_pattern_0 : IN STD_LOGIC;
    ctl_tx_test_pattern_1 : IN STD_LOGIC;
    ctl_tx_test_pattern_2 : IN STD_LOGIC;
    ctl_tx_test_pattern_3 : IN STD_LOGIC;
    ctl_tx_test_pattern_enable_0 : IN STD_LOGIC;
    ctl_tx_test_pattern_enable_1 : IN STD_LOGIC;
    ctl_tx_test_pattern_enable_2 : IN STD_LOGIC;
    ctl_tx_test_pattern_enable_3 : IN STD_LOGIC;
    ctl_tx_test_pattern_select_0 : IN STD_LOGIC;
    ctl_tx_test_pattern_select_1 : IN STD_LOGIC;
    ctl_tx_test_pattern_select_2 : IN STD_LOGIC;
    ctl_tx_test_pattern_select_3 : IN STD_LOGIC;
    ctl_tx_data_pattern_select_0 : IN STD_LOGIC;
    ctl_tx_data_pattern_select_1 : IN STD_LOGIC;
    ctl_tx_data_pattern_select_2 : IN STD_LOGIC;
    ctl_tx_data_pattern_select_3 : IN STD_LOGIC;
    ctl_tx_test_pattern_seed_a_0 : IN STD_LOGIC_VECTOR(57 DOWNTO 0);
    ctl_tx_test_pattern_seed_a_1 : IN STD_LOGIC_VECTOR(57 DOWNTO 0);
    ctl_tx_test_pattern_seed_a_2 : IN STD_LOGIC_VECTOR(57 DOWNTO 0);
    ctl_tx_test_pattern_seed_a_3 : IN STD_LOGIC_VECTOR(57 DOWNTO 0);
    ctl_tx_test_pattern_seed_b_0 : IN STD_LOGIC_VECTOR(57 DOWNTO 0);
    ctl_tx_test_pattern_seed_b_1 : IN STD_LOGIC_VECTOR(57 DOWNTO 0);
    ctl_tx_test_pattern_seed_b_2 : IN STD_LOGIC_VECTOR(57 DOWNTO 0);
    ctl_tx_test_pattern_seed_b_3 : IN STD_LOGIC_VECTOR(57 DOWNTO 0);
    ctl_tx_ipg_value_0 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    ctl_tx_ipg_value_1 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    ctl_tx_ipg_value_2 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    ctl_tx_ipg_value_3 : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    ctl_tx_custom_preamble_enable_0 : IN STD_LOGIC;
    ctl_tx_custom_preamble_enable_1 : IN STD_LOGIC;
    ctl_tx_custom_preamble_enable_2 : IN STD_LOGIC;
    ctl_tx_custom_preamble_enable_3 : IN STD_LOGIC;
    gt_loopback_in_0 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    gt_loopback_in_1 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    gt_loopback_in_2 : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    gt_loopback_in_3 : IN STD_LOGIC_VECTOR(2 DOWNTO 0)
  );
END COMPONENT;

END tech_mac_10g_quad_component_pkg;

