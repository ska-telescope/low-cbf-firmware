-------------------------------------------------------------------------------
-- Title      : CMAC Time division Multiplexing Package
-- Project    : 
-------------------------------------------------------------------------------
-- File       : cmac_tdm_pkg.vhd
-- Author     : William Kamp  <william.kamp@aut.ac.nz>
-- Company    : High Performance Computing Research Lab, Auckland University of Technology
-- Created    : 2017-05-05
-- Last update: 2018-05-18
-- Platform   : 
-- Standard   : VHDL'08
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Copyright (c) 2017 High Performance Computing Research Lab, Auckland University of Technology
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2017-05-05  1.0      will	Created
-- 2019-09-16  2.0p     nabel   Ported to Perentie
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.misc_tools_pkg.all;                  -- ceil_log2

package cmac_tdm_pkg is

    -- Package constants. Increase if required.
    constant pc_MAX_NUM_SAMPLES : natural := 128;
    constant pc_MAX_ANTENNA_PER_COL : natural := 10;

    type t_tdm_rd_ctrl is record
        rd_enable   : std_logic;
        dbl_buf_sel : std_logic;
        rd_addr     : unsigned(10 downto 0);  -- (ceil_log2(pc_MAX_ANTENNA_PER_COL*pc_MAX_NUM_SAMPLES)-1 downto 0);
        auto_corr   : std_logic;
        --pol_left    : std_logic;
        --pol_right   : std_logic;
        sample_cnt  : unsigned(7 downto 0);  -- (ceil_log2(pc_MAX_NUM_SAMPLES)-1 downto 0));
        sample_last : std_logic;
    end record t_tdm_rd_ctrl;
    
    type t_tdm_cache_wr_bus is record
        real_polX   : signed(8 downto 0);     -- (g_SAMPLE_WIDTH-1 downto 0);
        imag_polX   : signed(8 downto 0);     -- (g_SAMPLE_WIDTH-1 downto 0);
        real_polY   : signed(8 downto 0);     -- (g_SAMPLE_WIDTH-1 downto 0);
        imag_polY   : signed(8 downto 0);     -- (g_SAMPLE_WIDTH-1 downto 0);
        dbl_buf_sel : std_logic;
        wr_addr     : unsigned(15 downto 0);  -- (ceil_log2(g_NUM_SAMPLES*g_ANTENNA_PER_COL)-1 downto 0);
        wr_enable   : std_logic;
    end record t_tdm_cache_wr_bus;

    
    -- autogen start decl
 --------------------------------------------------
 -- Auto-generated code below. You should not edit.
 -- Generated Tue Aug  1 16:02:13 2017
 --------------------------------------------------
type t_tdm_rd_ctrl_a is array(natural range <>) of t_tdm_rd_ctrl;

constant T_TDM_RD_CTRL_ZERO : t_tdm_rd_ctrl := (
	rd_enable => '0',
	dbl_buf_sel => '0',
	rd_addr => (others => '0'),
	auto_corr => '0',
	sample_cnt => (others => '0'),
	sample_last => '0'
	);

constant T_TDM_RD_CTRL_SLV_WIDTH : natural := 23;

subtype t_tdm_rd_ctrl_slv is std_logic_vector(22 downto 0);
function to_slv (rec : t_tdm_rd_ctrl) return t_tdm_rd_ctrl_slv;

function from_slv (slv : std_logic_vector) return t_tdm_rd_ctrl;

type t_tdm_cache_wr_bus_a is array(natural range <>) of t_tdm_cache_wr_bus;

constant T_TDM_CACHE_WR_BUS_ZERO : t_tdm_cache_wr_bus := (
	real_polX => (others => '0'),
	imag_polX => (others => '0'),
	real_polY => (others => '0'),
	imag_polY => (others => '0'),
	dbl_buf_sel => '0',
	wr_addr => (others => '0'),
	wr_enable => '0'
	);

constant T_TDM_CACHE_WR_BUS_SLV_WIDTH : natural := 54;

subtype t_tdm_cache_wr_bus_slv is std_logic_vector(53 downto 0);
function to_slv (rec : t_tdm_cache_wr_bus) return t_tdm_cache_wr_bus_slv;

function from_slv (slv : std_logic_vector) return t_tdm_cache_wr_bus;

 ------------------------------------------------------
 -- End of Autogenerated code. You may add yours below.
 ------------------------------------------------------
    -- autogen end decl

    function f_ADDR_STRIDE (
        constant c_ANTENNA_PER_COL : natural;
        constant c_MAX_NUM_SAMPLES : natural)        
        return natural;
    
end package cmac_tdm_pkg;

package body cmac_tdm_pkg is

    -- autogen start body
 --------------------------------------------------
 -- Auto-generated code below. You should not edit.
 -- Generated Tue Aug  1 16:02:13 2017
 --------------------------------------------------
function to_slv (rec : t_tdm_rd_ctrl) return t_tdm_rd_ctrl_slv is
    variable slv : std_logic_vector(22 downto 0);
begin
    slv(0) := rec.sample_last;
    slv(8 downto 1) := std_logic_vector(rec.sample_cnt);
    slv(9) := rec.auto_corr;
    slv(20 downto 10) := std_logic_vector(rec.rd_addr);
    slv(21) := rec.dbl_buf_sel;
    slv(22) := rec.rd_enable;
return slv;
end function to_slv;

function from_slv (slv : std_logic_vector) return t_tdm_rd_ctrl is
    variable rec : t_tdm_rd_ctrl;
begin
    rec.sample_last := slv(0);
    rec.sample_cnt := unsigned(slv(8 downto 1));
    rec.auto_corr := slv(9);
    rec.rd_addr := unsigned(slv(20 downto 10));
    rec.dbl_buf_sel := slv(21);
    rec.rd_enable := slv(22);
return rec;
end function from_slv;

function to_slv (rec : t_tdm_cache_wr_bus) return t_tdm_cache_wr_bus_slv is
    variable slv : std_logic_vector(53 downto 0);
begin
    slv(0) := rec.wr_enable;
    slv(16 downto 1) := std_logic_vector(rec.wr_addr);
    slv(17) := rec.dbl_buf_sel;
    slv(26 downto 18) := std_logic_vector(rec.imag_polY);
    slv(35 downto 27) := std_logic_vector(rec.real_polY);
    slv(44 downto 36) := std_logic_vector(rec.imag_polX);
    slv(53 downto 45) := std_logic_vector(rec.real_polX);
return slv;
end function to_slv;

function from_slv (slv : std_logic_vector) return t_tdm_cache_wr_bus is
    variable rec : t_tdm_cache_wr_bus;
begin
    rec.wr_enable := slv(0);
    rec.wr_addr := unsigned(slv(16 downto 1));
    rec.dbl_buf_sel := slv(17);
    rec.imag_polY := signed(slv(26 downto 18));
    rec.real_polY := signed(slv(35 downto 27));
    rec.imag_polX := signed(slv(44 downto 36));
    rec.real_polX := signed(slv(53 downto 45));
return rec;
end function from_slv;

 ------------------------------------------------------
 -- End of Autogenerated code. You may add yours below.
 ------------------------------------------------------
    -- autogen end body

    function f_ADDR_STRIDE (
        constant c_ANTENNA_PER_COL : natural;
        constant c_MAX_NUM_SAMPLES : natural)        
        return natural is
    begin
        return 2**ceil_log2((c_ANTENNA_PER_COL-1)*c_MAX_NUM_SAMPLES)/(c_ANTENNA_PER_COL-1);
    end function;
    
end package body cmac_tdm_pkg;
