LIBRARY IEEE, technology_lib;
USE IEEE.std_logic_1164.ALL;
USE technology_lib.technology_pkg.ALL;


PACKAGE tech_mac_40g_pkg IS

   TYPE t_quad_locations_40g IS (
      QUAD_40G_122, QUAD_40G_124, QUAD_40G_125, QUAD_40G_126, QUAD_40G_128, QUAD_40G_130, QUAD_40G_131, QUAD_40G_132, QUAD_40G_134, QUAD_40G_135);


END tech_mac_40g_pkg;

