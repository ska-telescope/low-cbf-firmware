-------------------------------------------------------------
-- Ethernet CRC32 calculate and check 
-- Creation date 2019-07-12 23:39:50.054208
-- Written by python script : interconnectFCS.py
-- By David Humphrey (dave.humphrey@csiro.au) 
-- 
-- 
------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity crc32Full64Step is
   port (
      clk     : in std_logic;
      data_i  : in std_logic_vector(63 downto 0);
      valid_i : in std_logic;
      sof_i   : in std_logic;
      state_o : out std_logic_vector(31 downto 0);
      new_state_o : out std_logic_vector(31 downto 0) -- logic only path from data_i, bytes_i
   );
end crc32Full64Step;

architecture Behavioral of crc32Full64Step is

   signal allbits : std_logic_vector(95 downto 0);
   signal cur_state : std_logic_vector(31 downto 0);
   signal new_state : std_logic_vector(31 downto 0);
   signal LUT_gen0 : std_logic_vector(15 downto 0);
   signal LUT_gen0_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen0_block0_data : std_logic_vector(63 downto 0) := "1100110000110011001100111100110011001100001100110011001111001100";
   signal LUT_gen0_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen0_block1_data : std_logic_vector(63 downto 0) := "0101010110101010101010100101010110101010010101010101010110101010";
   signal LUT_gen0_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen0_block2_data : std_logic_vector(63 downto 0) := "1111000011110000000011110000111100001111000011111111000011110000";
   signal LUT_gen0_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen0_block3_data : std_logic_vector(63 downto 0) := "0011110000111100001111000011110000111100001111000011110000111100";
   signal LUT_gen0_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen0_block4_data : std_logic_vector(63 downto 0) := "1111111100000000111111110000000011111111000000001111111100000000";
   signal LUT_gen0_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen0_block5_data : std_logic_vector(63 downto 0) := "1010101001010101101010100101010101010101101010100101010110101010";
   signal LUT_gen0_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen0_block6_data : std_logic_vector(63 downto 0) := "1010010110100101101001011010010101011010010110100101101001011010";
   signal LUT_gen0_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen0_block7_data : std_logic_vector(63 downto 0) := "1001100110011001011001100110011010011001100110010110011001100110";
   signal LUT_gen0_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen0_block8_data : std_logic_vector(63 downto 0) := "0110011010011001100110010110011001100110100110011001100101100110";
   signal LUT_gen0_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen0_block9_data : std_logic_vector(63 downto 0) := "1111111111111111111111111111111100000000000000000000000000000000";
   signal LUT_gen0_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen0_block10_data : std_logic_vector(63 downto 0) := "1111000011110000000011110000111100001111000011111111000011110000";
   signal LUT_gen0_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen0_block11_data : std_logic_vector(63 downto 0) := "1001011010010110011010010110100101101001011010011001011010010110";
   signal LUT_gen0_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen0_block12_data : std_logic_vector(63 downto 0) := "1010101010101010101010101010101010101010101010101010101010101010";
   signal LUT_gen0_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen0_block13_data : std_logic_vector(63 downto 0) := "1111000011110000111100001111000011110000111100001111000011110000";
   signal LUT_gen0_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen0_block14_data : std_logic_vector(63 downto 0) := "1010010101011010101001010101101010100101010110101010010101011010";
   signal LUT_gen0_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen0_block15_data : std_logic_vector(63 downto 0) := "1010101010101010101010101010101010101010101010101010101010101010";
   signal LUT_gen1 : std_logic_vector(15 downto 0);
   signal LUT_gen1_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen1_block0_data : std_logic_vector(63 downto 0) := "0101101001011010101001011010010110100101101001010101101001011010";
   signal LUT_gen1_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen1_block1_data : std_logic_vector(63 downto 0) := "1100110011001100001100110011001100110011001100111100110011001100";
   signal LUT_gen1_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen1_block2_data : std_logic_vector(63 downto 0) := "1010101001010101101010100101010101010101101010100101010110101010";
   signal LUT_gen1_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen1_block3_data : std_logic_vector(63 downto 0) := "1010010101011010101001010101101010100101010110101010010101011010";
   signal LUT_gen1_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen1_block4_data : std_logic_vector(63 downto 0) := "1111111111111111000000000000000011111111111111110000000000000000";
   signal LUT_gen1_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen1_block5_data : std_logic_vector(63 downto 0) := "1100001111000011001111000011110011000011110000110011110000111100";
   signal LUT_gen1_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen1_block6_data : std_logic_vector(63 downto 0) := "1001100101100110100110010110011010011001011001101001100101100110";
   signal LUT_gen1_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen1_block7_data : std_logic_vector(63 downto 0) := "0110100101101001011010010110100110010110100101101001011010010110";
   signal LUT_gen1_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen1_block8_data : std_logic_vector(63 downto 0) := "0011110000111100110000111100001111000011110000110011110000111100";
   signal LUT_gen1_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen1_block10_data : std_logic_vector(63 downto 0) := "1010101001010101101010100101010101010101101010100101010110101010";
   signal LUT_gen1_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen1_block11_data : std_logic_vector(63 downto 0) := "1001011001101001100101100110100101101001100101100110100110010110";
   signal LUT_gen1_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen1_block12_data : std_logic_vector(63 downto 0) := "0110011001100110011001100110011001100110011001100110011001100110";
   signal LUT_gen1_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen1_block13_data : std_logic_vector(63 downto 0) := "1111111100000000111111110000000011111111000000001111111100000000";
   signal LUT_gen1_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen1_block14_data : std_logic_vector(63 downto 0) := "1100110000110011001100111100110011001100001100110011001111001100";
   signal LUT_gen1_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen1_block15_data : std_logic_vector(63 downto 0) := "1100110011001100110011001100110011001100110011001100110011001100";
   signal LUT_gen2 : std_logic_vector(15 downto 0);
   signal LUT_gen2_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen2_block0_data : std_logic_vector(63 downto 0) := "0110011010011001011001101001100110011001011001101001100101100110";
   signal LUT_gen2_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen2_block1_data : std_logic_vector(63 downto 0) := "1010010110100101101001011010010101011010010110100101101001011010";
   signal LUT_gen2_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen2_block2_data : std_logic_vector(63 downto 0) := "1001100110011001011001100110011010011001100110010110011001100110";
   signal LUT_gen2_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen2_block3_data : std_logic_vector(63 downto 0) := "0110011010011001100110010110011001100110100110011001100101100110";
   signal LUT_gen2_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen2_block4_data : std_logic_vector(63 downto 0) := "1111111111111111111111111111111100000000000000000000000000000000";
   signal LUT_gen2_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen2_block5_data : std_logic_vector(63 downto 0) := "1111000000001111111100000000111100001111111100000000111111110000";
   signal LUT_gen2_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen2_block6_data : std_logic_vector(63 downto 0) := "1100001111000011001111000011110011000011110000110011110000111100";
   signal LUT_gen2_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen2_block7_data : std_logic_vector(63 downto 0) := "1100001100111100110000110011110011000011001111001100001100111100";
   signal LUT_gen2_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen2_block8_data : std_logic_vector(63 downto 0) := "0101101010100101010110101010010110100101010110101010010101011010";
   signal LUT_gen2_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen2_block9_data : std_logic_vector(63 downto 0) := "1010101010101010101010101010101010101010101010101010101010101010";
   signal LUT_gen2_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen2_block10_data : std_logic_vector(63 downto 0) := "0011001100110011110011001100110000110011001100111100110011001100";
   signal LUT_gen2_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen2_block11_data : std_logic_vector(63 downto 0) := "1001011001101001011010011001011010010110011010010110100110010110";
   signal LUT_gen2_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen2_block12_data : std_logic_vector(63 downto 0) := "1001011010010110100101101001011010010110100101101001011010010110";
   signal LUT_gen2_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen2_block13_data : std_logic_vector(63 downto 0) := "1111111111111111000000000000000011111111111111110000000000000000";
   signal LUT_gen2_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen2_block14_data : std_logic_vector(63 downto 0) := "1111000011110000000011110000111100001111000011111111000011110000";
   signal LUT_gen2_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen2_block15_data : std_logic_vector(63 downto 0) := "1111000011110000111100001111000011110000111100001111000011110000";
   signal LUT_gen3 : std_logic_vector(15 downto 0);
   signal LUT_gen3_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen3_block0_data : std_logic_vector(63 downto 0) := "0110100101101001100101101001011001101001011010011001011010010110";
   signal LUT_gen3_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen3_block1_data : std_logic_vector(63 downto 0) := "1001100101100110100110010110011010011001011001101001100101100110";
   signal LUT_gen3_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen3_block2_data : std_logic_vector(63 downto 0) := "0110100101101001011010010110100110010110100101101001011010010110";
   signal LUT_gen3_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen3_block3_data : std_logic_vector(63 downto 0) := "0011110000111100110000111100001111000011110000110011110000111100";
   signal LUT_gen3_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen3_block5_data : std_logic_vector(63 downto 0) := "0101101010100101101001010101101001011010101001011010010101011010";
   signal LUT_gen3_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen3_block6_data : std_logic_vector(63 downto 0) := "0101101010100101010110101010010110100101010110101010010101011010";
   signal LUT_gen3_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen3_block7_data : std_logic_vector(63 downto 0) := "1111000000001111000011111111000011110000000011110000111111110000";
   signal LUT_gen3_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen3_block8_data : std_logic_vector(63 downto 0) := "1100110000110011001100111100110011001100001100110011001111001100";
   signal LUT_gen3_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen3_block9_data : std_logic_vector(63 downto 0) := "0110011001100110011001100110011001100110011001100110011001100110";
   signal LUT_gen3_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen3_block10_data : std_logic_vector(63 downto 0) := "0000111100001111000011110000111111110000111100001111000011110000";
   signal LUT_gen3_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen3_block11_data : std_logic_vector(63 downto 0) := "1100001100111100001111001100001100111100110000111100001100111100";
   signal LUT_gen3_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen3_block12_data : std_logic_vector(63 downto 0) := "1100001100111100110000110011110011000011001111001100001100111100";
   signal LUT_gen3_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen3_block13_data : std_logic_vector(63 downto 0) := "1111111111111111111111111111111100000000000000000000000000000000";
   signal LUT_gen3_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen3_block14_data : std_logic_vector(63 downto 0) := "0000000011111111000000001111111111111111000000001111111100000000";
   signal LUT_gen3_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen3_block15_data : std_logic_vector(63 downto 0) := "0101010110101010010101011010101001010101101010100101010110101010";
   signal LUT_gen4 : std_logic_vector(15 downto 0);
   signal LUT_gen4_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen4_block0_data : std_logic_vector(63 downto 0) := "1001011001101001100101100110100101101001100101100110100110010110";
   signal LUT_gen4_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen4_block1_data : std_logic_vector(63 downto 0) := "1100001111000011001111000011110011000011110000110011110000111100";
   signal LUT_gen4_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen4_block2_data : std_logic_vector(63 downto 0) := "1100001100111100110000110011110011000011001111001100001100111100";
   signal LUT_gen4_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen4_block3_data : std_logic_vector(63 downto 0) := "0101101010100101010110101010010110100101010110101010010101011010";
   signal LUT_gen4_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen4_block4_data : std_logic_vector(63 downto 0) := "1010101010101010101010101010101010101010101010101010101010101010";
   signal LUT_gen4_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen4_block5_data : std_logic_vector(63 downto 0) := "1100001100111100001111001100001100111100110000111100001100111100";
   signal LUT_gen4_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen4_block6_data : std_logic_vector(63 downto 0) := "1100110000110011001100111100110011001100001100110011001111001100";
   signal LUT_gen4_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen4_block7_data : std_logic_vector(63 downto 0) := "0101010110101010101010100101010110101010010101010101010110101010";
   signal LUT_gen4_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen4_block8_data : std_logic_vector(63 downto 0) := "1111000011110000000011110000111100001111000011111111000011110000";
   signal LUT_gen4_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen4_block9_data : std_logic_vector(63 downto 0) := "0011110000111100001111000011110000111100001111000011110000111100";
   signal LUT_gen4_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen4_block10_data : std_logic_vector(63 downto 0) := "1111111100000000111111110000000011111111000000001111111100000000";
   signal LUT_gen4_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen4_block11_data : std_logic_vector(63 downto 0) := "1010010101011010010110101010010101011010101001011010010101011010";
   signal LUT_gen4_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen4_block12_data : std_logic_vector(63 downto 0) := "0101101010100101101001010101101001011010101001011010010101011010";
   signal LUT_gen4_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen4_block14_data : std_logic_vector(63 downto 0) := "0101010101010101101010101010101001010101010101011010101010101010";
   signal LUT_gen4_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen4_block15_data : std_logic_vector(63 downto 0) := "1001100110011001011001100110011010011001100110010110011001100110";
   signal LUT_gen5 : std_logic_vector(15 downto 0);
   signal LUT_gen5_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen5_block0_data : std_logic_vector(63 downto 0) := "0011110011000011110000110011110000111100110000111100001100111100";
   signal LUT_gen5_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen5_block1_data : std_logic_vector(63 downto 0) := "0101101010100101010110101010010110100101010110101010010101011010";
   signal LUT_gen5_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen5_block2_data : std_logic_vector(63 downto 0) := "1111000000001111000011111111000011110000000011110000111111110000";
   signal LUT_gen5_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen5_block3_data : std_logic_vector(63 downto 0) := "1100110000110011001100111100110011001100001100110011001111001100";
   signal LUT_gen5_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen5_block4_data : std_logic_vector(63 downto 0) := "0110011001100110011001100110011001100110011001100110011001100110";
   signal LUT_gen5_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen5_block5_data : std_logic_vector(63 downto 0) := "1111111100000000000000001111111100000000111111111111111100000000";
   signal LUT_gen5_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen5_block6_data : std_logic_vector(63 downto 0) := "0101101001011010101001011010010110100101101001010101101001011010";
   signal LUT_gen5_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen5_block7_data : std_logic_vector(63 downto 0) := "1100110011001100001100110011001100110011001100111100110011001100";
   signal LUT_gen5_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen5_block8_data : std_logic_vector(63 downto 0) := "1010101001010101101010100101010101010101101010100101010110101010";
   signal LUT_gen5_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen5_block9_data : std_logic_vector(63 downto 0) := "1010010101011010101001010101101010100101010110101010010101011010";
   signal LUT_gen5_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen5_block10_data : std_logic_vector(63 downto 0) := "1111111111111111000000000000000011111111111111110000000000000000";
   signal LUT_gen5_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen5_block11_data : std_logic_vector(63 downto 0) := "0011001111001100110011000011001111001100001100110011001111001100";
   signal LUT_gen5_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen5_block12_data : std_logic_vector(63 downto 0) := "1001100101100110011001101001100101100110100110011001100101100110";
   signal LUT_gen5_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen5_block14_data : std_logic_vector(63 downto 0) := "0011001100110011001100110011001111001100110011001100110011001100";
   signal LUT_gen5_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen5_block15_data : std_logic_vector(63 downto 0) := "1100001111000011110000111100001100111100001111000011110000111100";
   signal LUT_gen6 : std_logic_vector(15 downto 0);
   signal LUT_gen6_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen6_block0_data : std_logic_vector(63 downto 0) := "1100001111000011110000111100001100111100001111000011110000111100";
   signal LUT_gen6_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen6_block1_data : std_logic_vector(63 downto 0) := "1001100110011001100110011001100101100110011001100110011001100110";
   signal LUT_gen6_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen6_block2_data : std_logic_vector(63 downto 0) := "1010010101011010101001010101101010100101010110101010010101011010";
   signal LUT_gen6_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen6_block3_data : std_logic_vector(63 downto 0) := "1100110011001100001100110011001100110011001100111100110011001100";
   signal LUT_gen6_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen6_block4_data : std_logic_vector(63 downto 0) := "1100001100111100110000110011110011000011001111001100001100111100";
   signal LUT_gen6_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen6_block5_data : std_logic_vector(63 downto 0) := "1010101001010101010101011010101010101010010101010101010110101010";
   signal LUT_gen6_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen6_block6_data : std_logic_vector(63 downto 0) := "1100001100111100110000110011110011000011001111001100001100111100";
   signal LUT_gen6_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen6_block7_data : std_logic_vector(63 downto 0) := "0011110000111100110000111100001111000011110000110011110000111100";
   signal LUT_gen6_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen6_block8_data : std_logic_vector(63 downto 0) := "1111111100000000111111110000000011111111000000001111111100000000";
   signal LUT_gen6_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen6_block9_data : std_logic_vector(63 downto 0) := "1001100101100110011001101001100101100110100110011001100101100110";
   signal LUT_gen6_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen6_block10_data : std_logic_vector(63 downto 0) := "0000111100001111111100001111000000001111000011111111000011110000";
   signal LUT_gen6_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen6_block11_data : std_logic_vector(63 downto 0) := "0110011001100110011001100110011001100110011001100110011001100110";
   signal LUT_gen6_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen6_block12_data : std_logic_vector(63 downto 0) := "0011110000111100110000111100001111000011110000110011110000111100";
   signal LUT_gen6_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen6_block13_data : std_logic_vector(63 downto 0) := "0101101001011010010110100101101001011010010110100101101001011010";
   signal LUT_gen6_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen6_block14_data : std_logic_vector(63 downto 0) := "0101010110101010010101011010101001010101101010100101010110101010";
   signal LUT_gen6_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen6_block15_data : std_logic_vector(63 downto 0) := "0000111111110000000011111111000000001111111100000000111111110000";
   signal LUT_gen7 : std_logic_vector(15 downto 0);
   signal LUT_gen7_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen7_block0_data : std_logic_vector(63 downto 0) := "1010010101011010101001010101101010100101010110101010010101011010";
   signal LUT_gen7_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen7_block1_data : std_logic_vector(63 downto 0) := "1001011010010110100101101001011010010110100101101001011010010110";
   signal LUT_gen7_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen7_block2_data : std_logic_vector(63 downto 0) := "0110011010011001100110010110011001100110100110011001100101100110";
   signal LUT_gen7_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen7_block3_data : std_logic_vector(63 downto 0) := "0000111100001111000011110000111111110000111100001111000011110000";
   signal LUT_gen7_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen7_block4_data : std_logic_vector(63 downto 0) := "0101101010100101101001010101101001011010101001011010010101011010";
   signal LUT_gen7_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen7_block5_data : std_logic_vector(63 downto 0) := "0011110000111100110000111100001111000011110000110011110000111100";
   signal LUT_gen7_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen7_block6_data : std_logic_vector(63 downto 0) := "1111000000001111000011111111000011110000000011110000111111110000";
   signal LUT_gen7_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen7_block7_data : std_logic_vector(63 downto 0) := "1111000000001111111100000000111100001111111100000000111111110000";
   signal LUT_gen7_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen7_block8_data : std_logic_vector(63 downto 0) := "0101010101010101101010101010101001010101010101011010101010101010";
   signal LUT_gen7_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen7_block9_data : std_logic_vector(63 downto 0) := "0011110000111100110000111100001111000011110000110011110000111100";
   signal LUT_gen7_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen7_block10_data : std_logic_vector(63 downto 0) := "1010101001010101101010100101010101010101101010100101010110101010";
   signal LUT_gen7_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen7_block11_data : std_logic_vector(63 downto 0) := "0011110000111100001111000011110000111100001111000011110000111100";
   signal LUT_gen7_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen7_block12_data : std_logic_vector(63 downto 0) := "1111000000001111111100000000111100001111111100000000111111110000";
   signal LUT_gen7_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen7_block13_data : std_logic_vector(63 downto 0) := "1001100101100110100110010110011010011001011001101001100101100110";
   signal LUT_gen7_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen7_block14_data : std_logic_vector(63 downto 0) := "0011001100110011110011001100110000110011001100111100110011001100";
   signal LUT_gen7_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen7_block15_data : std_logic_vector(63 downto 0) := "0000000011111111111111110000000000000000111111111111111100000000";
   signal LUT_gen8 : std_logic_vector(15 downto 0);
   signal LUT_gen8_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen8_block0_data : std_logic_vector(63 downto 0) := "1100110000110011001100111100110011001100001100110011001111001100";
   signal LUT_gen8_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen8_block1_data : std_logic_vector(63 downto 0) := "1100001100111100110000110011110011000011001111001100001100111100";
   signal LUT_gen8_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen8_block2_data : std_logic_vector(63 downto 0) := "0011110000111100110000111100001111000011110000110011110000111100";
   signal LUT_gen8_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen8_block3_data : std_logic_vector(63 downto 0) := "1111111100000000111111110000000011111111000000001111111100000000";
   signal LUT_gen8_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen8_block4_data : std_logic_vector(63 downto 0) := "1001100101100110011001101001100101100110100110011001100101100110";
   signal LUT_gen8_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen8_block5_data : std_logic_vector(63 downto 0) := "0000000011111111000000001111111111111111000000001111111100000000";
   signal LUT_gen8_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen8_block6_data : std_logic_vector(63 downto 0) := "0101010110101010101010100101010110101010010101010101010110101010";
   signal LUT_gen8_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen8_block7_data : std_logic_vector(63 downto 0) := "0000000011111111111111110000000000000000111111111111111100000000";
   signal LUT_gen8_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen8_block8_data : std_logic_vector(63 downto 0) := "1001100110011001100110011001100101100110011001100110011001100110";
   signal LUT_gen8_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen8_block9_data : std_logic_vector(63 downto 0) := "1111000000001111111100000000111100001111111100000000111111110000";
   signal LUT_gen8_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen8_block10_data : std_logic_vector(63 downto 0) := "1001100110011001011001100110011010011001100110010110011001100110";
   signal LUT_gen8_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen8_block11_data : std_logic_vector(63 downto 0) := "1010010101011010101001010101101010100101010110101010010101011010";
   signal LUT_gen8_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen8_block12_data : std_logic_vector(63 downto 0) := "0000000011111111111111110000000000000000111111111111111100000000";
   signal LUT_gen8_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen8_block13_data : std_logic_vector(63 downto 0) := "0110100101101001100101101001011001101001011010011001011010010110";
   signal LUT_gen8_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen8_block14_data : std_logic_vector(63 downto 0) := "0000111100001111000011110000111111110000111100001111000011110000";
   signal LUT_gen8_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen8_block15_data : std_logic_vector(63 downto 0) := "0000000000000000111111111111111111111111111111110000000000000000";
   signal LUT_gen9 : std_logic_vector(15 downto 0);
   signal LUT_gen9_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen9_block0_data : std_logic_vector(63 downto 0) := "0011110011000011001111001100001111000011001111001100001100111100";
   signal LUT_gen9_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen9_block1_data : std_logic_vector(63 downto 0) := "1010010110100101101001011010010101011010010110100101101001011010";
   signal LUT_gen9_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen9_block2_data : std_logic_vector(63 downto 0) := "0000000011111111111111110000000000000000111111111111111100000000";
   signal LUT_gen9_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen9_block3_data : std_logic_vector(63 downto 0) := "0110100101101001100101101001011001101001011010011001011010010110";
   signal LUT_gen9_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen9_block4_data : std_logic_vector(63 downto 0) := "1100001100111100001111001100001100111100110000111100001100111100";
   signal LUT_gen9_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen9_block5_data : std_logic_vector(63 downto 0) := "1111111100000000000000001111111100000000111111111111111100000000";
   signal LUT_gen9_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen9_block6_data : std_logic_vector(63 downto 0) := "1100001111000011001111000011110011000011110000110011110000111100";
   signal LUT_gen9_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen9_block7_data : std_logic_vector(63 downto 0) := "0011001100110011001100110011001111001100110011001100110011001100";
   signal LUT_gen9_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen9_block8_data : std_logic_vector(63 downto 0) := "0101101010100101101001010101101001011010101001011010010101011010";
   signal LUT_gen9_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen9_block9_data : std_logic_vector(63 downto 0) := "0101010110101010101010100101010110101010010101010101010110101010";
   signal LUT_gen9_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen9_block10_data : std_logic_vector(63 downto 0) := "1001100110011001011001100110011010011001100110010110011001100110";
   signal LUT_gen9_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen9_block11_data : std_logic_vector(63 downto 0) := "0101101010100101010110101010010110100101010110101010010101011010";
   signal LUT_gen9_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen9_block12_data : std_logic_vector(63 downto 0) := "1010101010101010010101010101010101010101010101011010101010101010";
   signal LUT_gen9_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen9_block13_data : std_logic_vector(63 downto 0) := "1100110000110011110011000011001100110011110011000011001111001100";
   signal LUT_gen9_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen9_block14_data : std_logic_vector(63 downto 0) := "0101101001011010010110100101101001011010010110100101101001011010";
   signal LUT_gen9_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen9_block15_data : std_logic_vector(63 downto 0) := "1111111111111111111111111111111100000000000000000000000000000000";
   signal LUT_gen10 : std_logic_vector(15 downto 0);
   signal LUT_gen10_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen10_block0_data : std_logic_vector(63 downto 0) := "0011110000111100001111000011110000111100001111000011110000111100";
   signal LUT_gen10_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen10_block1_data : std_logic_vector(63 downto 0) := "1100110011001100001100110011001100110011001100111100110011001100";
   signal LUT_gen10_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen10_block2_data : std_logic_vector(63 downto 0) := "0101101001011010010110100101101001011010010110100101101001011010";
   signal LUT_gen10_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen10_block3_data : std_logic_vector(63 downto 0) := "0000000011111111000000001111111111111111000000001111111100000000";
   signal LUT_gen10_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen10_block4_data : std_logic_vector(63 downto 0) := "1111000011110000000011110000111100001111000011111111000011110000";
   signal LUT_gen10_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen10_block5_data : std_logic_vector(63 downto 0) := "0000000011111111111111110000000000000000111111111111111100000000";
   signal LUT_gen10_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen10_block6_data : std_logic_vector(63 downto 0) := "1111111100000000111111110000000011111111000000001111111100000000";
   signal LUT_gen10_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen10_block7_data : std_logic_vector(63 downto 0) := "0110100101101001100101101001011001101001011010011001011010010110";
   signal LUT_gen10_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen10_block8_data : std_logic_vector(63 downto 0) := "1111111111111111111111111111111100000000000000000000000000000000";
   signal LUT_gen10_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen10_block9_data : std_logic_vector(63 downto 0) := "0011001100110011110011001100110000110011001100111100110011001100";
   signal LUT_gen10_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen10_block10_data : std_logic_vector(63 downto 0) := "1001100110011001011001100110011010011001100110010110011001100110";
   signal LUT_gen10_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen10_block11_data : std_logic_vector(63 downto 0) := "0101101010100101010110101010010110100101010110101010010101011010";
   signal LUT_gen10_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen10_block12_data : std_logic_vector(63 downto 0) := "0011001100110011001100110011001111001100110011001100110011001100";
   signal LUT_gen10_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen10_block13_data : std_logic_vector(63 downto 0) := "0101010101010101101010101010101001010101010101011010101010101010";
   signal LUT_gen10_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen10_block14_data : std_logic_vector(63 downto 0) := "0011110000111100001111000011110000111100001111000011110000111100";
   signal LUT_gen10_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen10_block15_data : std_logic_vector(63 downto 0) := "1010101010101010101010101010101010101010101010101010101010101010";
   signal LUT_gen11 : std_logic_vector(15 downto 0);
   signal LUT_gen11_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen11_block0_data : std_logic_vector(63 downto 0) := "0000111111110000000011111111000000001111111100000000111111110000";
   signal LUT_gen11_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen11_block1_data : std_logic_vector(63 downto 0) := "0000111100001111000011110000111111110000111100001111000011110000";
   signal LUT_gen11_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen11_block2_data : std_logic_vector(63 downto 0) := "1001100101100110100110010110011010011001011001101001100101100110";
   signal LUT_gen11_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen11_block3_data : std_logic_vector(63 downto 0) := "1111111111111111000000000000000011111111111111110000000000000000";
   signal LUT_gen11_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen11_block4_data : std_logic_vector(63 downto 0) := "1010101001010101101010100101010101010101101010100101010110101010";
   signal LUT_gen11_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen11_block5_data : std_logic_vector(63 downto 0) := "1010101010101010010101010101010101010101010101011010101010101010";
   signal LUT_gen11_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen11_block6_data : std_logic_vector(63 downto 0) := "1111111111111111000000000000000011111111111111110000000000000000";
   signal LUT_gen11_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen11_block7_data : std_logic_vector(63 downto 0) := "0011110011000011001111001100001111000011001111001100001100111100";
   signal LUT_gen11_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen11_block9_data : std_logic_vector(63 downto 0) := "1010010110100101101001011010010101011010010110100101101001011010";
   signal LUT_gen11_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen11_block10_data : std_logic_vector(63 downto 0) := "1100001111000011110000111100001100111100001111000011110000111100";
   signal LUT_gen11_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen11_block11_data : std_logic_vector(63 downto 0) := "1100110000110011001100111100110011001100001100110011001111001100";
   signal LUT_gen11_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen11_block12_data : std_logic_vector(63 downto 0) := "0101101001011010010110100101101001011010010110100101101001011010";
   signal LUT_gen11_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen11_block13_data : std_logic_vector(63 downto 0) := "1001100110011001100110011001100101100110011001100110011001100110";
   signal LUT_gen11_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen11_block14_data : std_logic_vector(63 downto 0) := "0000111111110000000011111111000000001111111100000000111111110000";
   signal LUT_gen11_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen11_block15_data : std_logic_vector(63 downto 0) := "1100110011001100110011001100110011001100110011001100110011001100";
   signal LUT_gen12 : std_logic_vector(15 downto 0);
   signal LUT_gen12_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen12_block0_data : std_logic_vector(63 downto 0) := "0000000011111111111111110000000000000000111111111111111100000000";
   signal LUT_gen12_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen12_block1_data : std_logic_vector(63 downto 0) := "1111111100000000111111110000000011111111000000001111111100000000";
   signal LUT_gen12_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen12_block2_data : std_logic_vector(63 downto 0) := "0110100101101001100101101001011001101001011010011001011010010110";
   signal LUT_gen12_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen12_block3_data : std_logic_vector(63 downto 0) := "1111111111111111111111111111111100000000000000000000000000000000";
   signal LUT_gen12_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen12_block4_data : std_logic_vector(63 downto 0) := "0011001100110011110011001100110000110011001100111100110011001100";
   signal LUT_gen12_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen12_block5_data : std_logic_vector(63 downto 0) := "1001100110011001100110011001100101100110011001100110011001100110";
   signal LUT_gen12_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen12_block6_data : std_logic_vector(63 downto 0) := "0101010101010101010101010101010110101010101010101010101010101010";
   signal LUT_gen12_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen12_block7_data : std_logic_vector(63 downto 0) := "1111000000001111000011111111000011110000000011110000111111110000";
   signal LUT_gen12_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen12_block8_data : std_logic_vector(63 downto 0) := "1010101010101010101010101010101010101010101010101010101010101010";
   signal LUT_gen12_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen12_block9_data : std_logic_vector(63 downto 0) := "0011001111001100001100111100110000110011110011000011001111001100";
   signal LUT_gen12_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen12_block10_data : std_logic_vector(63 downto 0) := "1010010101011010101001010101101010100101010110101010010101011010";
   signal LUT_gen12_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen12_block11_data : std_logic_vector(63 downto 0) := "0101101001011010101001011010010110100101101001010101101001011010";
   signal LUT_gen12_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen12_block12_data : std_logic_vector(63 downto 0) := "0011001111001100001100111100110000110011110011000011001111001100";
   signal LUT_gen12_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen12_block13_data : std_logic_vector(63 downto 0) := "0011110000111100001111000011110000111100001111000011110000111100";
   signal LUT_gen12_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen12_block14_data : std_logic_vector(63 downto 0) := "1010101001010101010101011010101010101010010101010101010110101010";
   signal LUT_gen12_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen12_block15_data : std_logic_vector(63 downto 0) := "1111000011110000111100001111000011110000111100001111000011110000";
   signal LUT_gen13 : std_logic_vector(15 downto 0);
   signal LUT_gen13_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen13_block0_data : std_logic_vector(63 downto 0) := "0000000000000000111111111111111111111111111111110000000000000000";
   signal LUT_gen13_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen13_block1_data : std_logic_vector(63 downto 0) := "1111111111111111000000000000000011111111111111110000000000000000";
   signal LUT_gen13_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen13_block2_data : std_logic_vector(63 downto 0) := "0011110011000011001111001100001111000011001111001100001100111100";
   signal LUT_gen13_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen13_block4_data : std_logic_vector(63 downto 0) := "1010010110100101101001011010010101011010010110100101101001011010";
   signal LUT_gen13_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen13_block5_data : std_logic_vector(63 downto 0) := "1100110011001100110011001100110011001100110011001100110011001100";
   signal LUT_gen13_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen13_block6_data : std_logic_vector(63 downto 0) := "0110011001100110011001100110011001100110011001100110011001100110";
   signal LUT_gen13_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen13_block7_data : std_logic_vector(63 downto 0) := "0101010110101010101010100101010110101010010101010101010110101010";
   signal LUT_gen13_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen13_block8_data : std_logic_vector(63 downto 0) := "1100110011001100110011001100110011001100110011001100110011001100";
   signal LUT_gen13_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen13_block9_data : std_logic_vector(63 downto 0) := "0000111100001111111100001111000000001111000011111111000011110000";
   signal LUT_gen13_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen13_block10_data : std_logic_vector(63 downto 0) := "1100110000110011001100111100110011001100001100110011001111001100";
   signal LUT_gen13_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen13_block11_data : std_logic_vector(63 downto 0) := "1100110000110011110011000011001100110011110011000011001111001100";
   signal LUT_gen13_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen13_block12_data : std_logic_vector(63 downto 0) := "1010010110100101010110100101101010100101101001010101101001011010";
   signal LUT_gen13_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen13_block13_data : std_logic_vector(63 downto 0) := "0000111111110000000011111111000000001111111100000000111111110000";
   signal LUT_gen13_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen13_block14_data : std_logic_vector(63 downto 0) := "1100110011001100001100110011001100110011001100111100110011001100";
   signal LUT_gen13_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen13_block15_data : std_logic_vector(63 downto 0) := "1111111100000000111111110000000011111111000000001111111100000000";
   signal LUT_gen14 : std_logic_vector(15 downto 0);
   signal LUT_gen14_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen14_block0_data : std_logic_vector(63 downto 0) := "1111111111111111111111111111111100000000000000000000000000000000";
   signal LUT_gen14_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen14_block1_data : std_logic_vector(63 downto 0) := "0101010101010101010101010101010110101010101010101010101010101010";
   signal LUT_gen14_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen14_block2_data : std_logic_vector(63 downto 0) := "1111000000001111000011111111000011110000000011110000111111110000";
   signal LUT_gen14_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen14_block3_data : std_logic_vector(63 downto 0) := "1010101010101010101010101010101010101010101010101010101010101010";
   signal LUT_gen14_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen14_block4_data : std_logic_vector(63 downto 0) := "0011001111001100001100111100110000110011110011000011001111001100";
   signal LUT_gen14_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen14_block5_data : std_logic_vector(63 downto 0) := "1010101010101010101010101010101010101010101010101010101010101010";
   signal LUT_gen14_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen14_block6_data : std_logic_vector(63 downto 0) := "0011110000111100001111000011110000111100001111000011110000111100";
   signal LUT_gen14_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen14_block7_data : std_logic_vector(63 downto 0) := "1100110011001100001100110011001100110011001100111100110011001100";
   signal LUT_gen14_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen14_block8_data : std_logic_vector(63 downto 0) := "0101101001011010010110100101101001011010010110100101101001011010";
   signal LUT_gen14_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen14_block9_data : std_logic_vector(63 downto 0) := "0000000011111111000000001111111111111111000000001111111100000000";
   signal LUT_gen14_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen14_block10_data : std_logic_vector(63 downto 0) := "1111000011110000000011110000111100001111000011111111000011110000";
   signal LUT_gen14_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen14_block11_data : std_logic_vector(63 downto 0) := "0000111100001111111100001111000000001111000011111111000011110000";
   signal LUT_gen14_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen14_block12_data : std_logic_vector(63 downto 0) := "0110011010011001011001101001100110011001011001101001100101100110";
   signal LUT_gen14_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen14_block13_data : std_logic_vector(63 downto 0) := "0000000011111111111111110000000000000000111111111111111100000000";
   signal LUT_gen14_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen14_block14_data : std_logic_vector(63 downto 0) := "0000111100001111000011110000111111110000111100001111000011110000";
   signal LUT_gen14_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen14_block15_data : std_logic_vector(63 downto 0) := "0101010101010101101010101010101001010101010101011010101010101010";
   signal LUT_gen15 : std_logic_vector(15 downto 0);
   signal LUT_gen15_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen15_block1_data : std_logic_vector(63 downto 0) := "0110011001100110011001100110011001100110011001100110011001100110";
   signal LUT_gen15_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen15_block2_data : std_logic_vector(63 downto 0) := "0101010110101010101010100101010110101010010101010101010110101010";
   signal LUT_gen15_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen15_block3_data : std_logic_vector(63 downto 0) := "1100110011001100110011001100110011001100110011001100110011001100";
   signal LUT_gen15_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen15_block4_data : std_logic_vector(63 downto 0) := "0000111100001111111100001111000000001111000011111111000011110000";
   signal LUT_gen15_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen15_block5_data : std_logic_vector(63 downto 0) := "1100110011001100110011001100110011001100110011001100110011001100";
   signal LUT_gen15_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen15_block6_data : std_logic_vector(63 downto 0) := "0000111111110000000011111111000000001111111100000000111111110000";
   signal LUT_gen15_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen15_block7_data : std_logic_vector(63 downto 0) := "0000111100001111000011110000111111110000111100001111000011110000";
   signal LUT_gen15_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen15_block8_data : std_logic_vector(63 downto 0) := "1001100101100110100110010110011010011001011001101001100101100110";
   signal LUT_gen15_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen15_block9_data : std_logic_vector(63 downto 0) := "1111111111111111000000000000000011111111111111110000000000000000";
   signal LUT_gen15_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen15_block10_data : std_logic_vector(63 downto 0) := "1010101001010101101010100101010101010101101010100101010110101010";
   signal LUT_gen15_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen15_block11_data : std_logic_vector(63 downto 0) := "1010101001010101101010100101010101010101101010100101010110101010";
   signal LUT_gen15_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen15_block12_data : std_logic_vector(63 downto 0) := "1100001111000011001111000011110011000011110000110011110000111100";
   signal LUT_gen15_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen15_block13_data : std_logic_vector(63 downto 0) := "1010101010101010010101010101010101010101010101011010101010101010";
   signal LUT_gen15_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen15_block14_data : std_logic_vector(63 downto 0) := "1111111100000000111111110000000011111111000000001111111100000000";
   signal LUT_gen15_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen15_block15_data : std_logic_vector(63 downto 0) := "1001100110011001100110011001100101100110011001100110011001100110";
   signal LUT_gen16 : std_logic_vector(15 downto 0);
   signal LUT_gen16_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen16_block0_data : std_logic_vector(63 downto 0) := "1100110000110011001100111100110011001100001100110011001111001100";
   signal LUT_gen16_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen16_block1_data : std_logic_vector(63 downto 0) := "0110100110010110100101100110100110010110011010010110100110010110";
   signal LUT_gen16_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen16_block2_data : std_logic_vector(63 downto 0) := "0011110000111100001111000011110000111100001111000011110000111100";
   signal LUT_gen16_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen16_block3_data : std_logic_vector(63 downto 0) := "0110011001100110011001100110011001100110011001100110011001100110";
   signal LUT_gen16_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen16_block4_data : std_logic_vector(63 downto 0) := "1111111111111111111111111111111100000000000000000000000000000000";
   signal LUT_gen16_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen16_block5_data : std_logic_vector(63 downto 0) := "1010101001010101101010100101010101010101101010100101010110101010";
   signal LUT_gen16_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen16_block6_data : std_logic_vector(63 downto 0) := "1010010101011010010110101010010101011010101001011010010101011010";
   signal LUT_gen16_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen16_block7_data : std_logic_vector(63 downto 0) := "0110011010011001100110010110011001100110100110011001100101100110";
   signal LUT_gen16_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen16_block8_data : std_logic_vector(63 downto 0) := "0000111111110000000011111111000000001111111100000000111111110000";
   signal LUT_gen16_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen16_block10_data : std_logic_vector(63 downto 0) := "1100001111000011110000111100001100111100001111000011110000111100";
   signal LUT_gen16_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen16_block11_data : std_logic_vector(63 downto 0) := "0000111100001111000011110000111111110000111100001111000011110000";
   signal LUT_gen16_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen16_block12_data : std_logic_vector(63 downto 0) := "1111000000001111111100000000111100001111111100000000111111110000";
   signal LUT_gen16_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen16_block13_data : std_logic_vector(63 downto 0) := "1100001111000011110000111100001100111100001111000011110000111100";
   signal LUT_gen16_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen16_block14_data : std_logic_vector(63 downto 0) := "1111000000001111000011111111000011110000000011110000111111110000";
   signal LUT_gen16_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen16_block15_data : std_logic_vector(63 downto 0) := "1001011010010110100101101001011010010110100101101001011010010110";
   signal LUT_gen17 : std_logic_vector(15 downto 0);
   signal LUT_gen17_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen17_block0_data : std_logic_vector(63 downto 0) := "0101101001011010101001011010010110100101101001010101101001011010";
   signal LUT_gen17_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen17_block1_data : std_logic_vector(63 downto 0) := "1100001100111100001111001100001100111100110000111100001100111100";
   signal LUT_gen17_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen17_block2_data : std_logic_vector(63 downto 0) := "1010010101011010101001010101101010100101010110101010010101011010";
   signal LUT_gen17_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen17_block3_data : std_logic_vector(63 downto 0) := "0011110000111100001111000011110000111100001111000011110000111100";
   signal LUT_gen17_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen17_block5_data : std_logic_vector(63 downto 0) := "0110100101101001100101101001011001101001011010011001011010010110";
   signal LUT_gen17_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen17_block6_data : std_logic_vector(63 downto 0) := "1001100101100110011001101001100101100110100110011001100101100110";
   signal LUT_gen17_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen17_block7_data : std_logic_vector(63 downto 0) := "1001011010010110011010010110100101101001011010011001011010010110";
   signal LUT_gen17_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen17_block8_data : std_logic_vector(63 downto 0) := "0000000011111111111111110000000000000000111111111111111100000000";
   signal LUT_gen17_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen17_block10_data : std_logic_vector(63 downto 0) := "0000111111110000000011111111000000001111111100000000111111110000";
   signal LUT_gen17_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen17_block11_data : std_logic_vector(63 downto 0) := "0101010110101010010101011010101001010101101010100101010110101010";
   signal LUT_gen17_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen17_block12_data : std_logic_vector(63 downto 0) := "1010101001010101010101011010101010101010010101010101010110101010";
   signal LUT_gen17_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen17_block13_data : std_logic_vector(63 downto 0) := "1010010101011010101001010101101010100101010110101010010101011010";
   signal LUT_gen17_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen17_block14_data : std_logic_vector(63 downto 0) := "0101010110101010101010100101010110101010010101010101010110101010";
   signal LUT_gen17_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen17_block15_data : std_logic_vector(63 downto 0) := "1100001100111100110000110011110011000011001111001100001100111100";
   signal LUT_gen18 : std_logic_vector(15 downto 0);
   signal LUT_gen18_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen18_block0_data : std_logic_vector(63 downto 0) := "1100110000110011110011000011001100110011110011000011001111001100";
   signal LUT_gen18_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen18_block1_data : std_logic_vector(63 downto 0) := "1010010101011010010110101010010101011010101001011010010101011010";
   signal LUT_gen18_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen18_block2_data : std_logic_vector(63 downto 0) := "0110011010011001100110010110011001100110100110011001100101100110";
   signal LUT_gen18_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen18_block3_data : std_logic_vector(63 downto 0) := "0000111111110000000011111111000000001111111100000000111111110000";
   signal LUT_gen18_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen18_block5_data : std_logic_vector(63 downto 0) := "1100110000110011110011000011001100110011110011000011001111001100";
   signal LUT_gen18_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen18_block6_data : std_logic_vector(63 downto 0) := "0011110000111100110000111100001111000011110000110011110000111100";
   signal LUT_gen18_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen18_block7_data : std_logic_vector(63 downto 0) := "1001011001101001100101100110100101101001100101100110100110010110";
   signal LUT_gen18_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen18_block8_data : std_logic_vector(63 downto 0) := "1010101010101010010101010101010101010101010101011010101010101010";
   signal LUT_gen18_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen18_block10_data : std_logic_vector(63 downto 0) := "0000000011111111111111110000000000000000111111111111111100000000";
   signal LUT_gen18_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen18_block11_data : std_logic_vector(63 downto 0) := "0011001100110011110011001100110000110011001100111100110011001100";
   signal LUT_gen18_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen18_block12_data : std_logic_vector(63 downto 0) := "1100110011001100001100110011001100110011001100111100110011001100";
   signal LUT_gen18_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen18_block13_data : std_logic_vector(63 downto 0) := "1100110000110011001100111100110011001100001100110011001111001100";
   signal LUT_gen18_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen18_block14_data : std_logic_vector(63 downto 0) := "1100110011001100001100110011001100110011001100111100110011001100";
   signal LUT_gen18_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen18_block15_data : std_logic_vector(63 downto 0) := "0101101010100101101001010101101001011010101001011010010101011010";
   signal LUT_gen19 : std_logic_vector(15 downto 0);
   signal LUT_gen19_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen19_block0_data : std_logic_vector(63 downto 0) := "1010010110100101010110100101101010100101101001010101101001011010";
   signal LUT_gen19_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen19_block1_data : std_logic_vector(63 downto 0) := "1001100101100110011001101001100101100110100110011001100101100110";
   signal LUT_gen19_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen19_block2_data : std_logic_vector(63 downto 0) := "1001011010010110011010010110100101101001011010011001011010010110";
   signal LUT_gen19_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen19_block3_data : std_logic_vector(63 downto 0) := "0000000011111111111111110000000000000000111111111111111100000000";
   signal LUT_gen19_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen19_block5_data : std_logic_vector(63 downto 0) := "0000111100001111111100001111000000001111000011111111000011110000";
   signal LUT_gen19_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen19_block6_data : std_logic_vector(63 downto 0) := "0101101010100101010110101010010110100101010110101010010101011010";
   signal LUT_gen19_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen19_block7_data : std_logic_vector(63 downto 0) := "1001011001101001011010011001011010010110011010010110100110010110";
   signal LUT_gen19_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen19_block8_data : std_logic_vector(63 downto 0) := "1001100110011001100110011001100101100110011001100110011001100110";
   signal LUT_gen19_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen19_block9_data : std_logic_vector(63 downto 0) := "1010101010101010101010101010101010101010101010101010101010101010";
   signal LUT_gen19_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen19_block10_data : std_logic_vector(63 downto 0) := "0000000000000000111111111111111111111111111111110000000000000000";
   signal LUT_gen19_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen19_block11_data : std_logic_vector(63 downto 0) := "0000111100001111000011110000111111110000111100001111000011110000";
   signal LUT_gen19_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen19_block12_data : std_logic_vector(63 downto 0) := "0000111100001111000011110000111111110000111100001111000011110000";
   signal LUT_gen19_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen19_block13_data : std_logic_vector(63 downto 0) := "0101101001011010101001011010010110100101101001010101101001011010";
   signal LUT_gen19_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen19_block14_data : std_logic_vector(63 downto 0) := "0000111100001111000011110000111111110000111100001111000011110000";
   signal LUT_gen19_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen19_block15_data : std_logic_vector(63 downto 0) := "1001100101100110011001101001100101100110100110011001100101100110";
   signal LUT_gen20 : std_logic_vector(15 downto 0);
   signal LUT_gen20_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen20_block0_data : std_logic_vector(63 downto 0) := "0000000000000000111111111111111111111111111111110000000000000000";
   signal LUT_gen20_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen20_block1_data : std_logic_vector(63 downto 0) := "0110100110010110011010011001011001101001100101100110100110010110";
   signal LUT_gen20_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen20_block2_data : std_logic_vector(63 downto 0) := "0110011010011001100110010110011001100110100110011001100101100110";
   signal LUT_gen20_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen20_block3_data : std_logic_vector(63 downto 0) := "1001011010010110011010010110100101101001011010011001011010010110";
   signal LUT_gen20_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen20_block4_data : std_logic_vector(63 downto 0) := "1111111100000000111111110000000011111111000000001111111100000000";
   signal LUT_gen20_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen20_block5_data : std_logic_vector(63 downto 0) := "1010101010101010101010101010101010101010101010101010101010101010";
   signal LUT_gen20_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen20_block6_data : std_logic_vector(63 downto 0) := "0110100110010110100101100110100110010110011010010110100110010110";
   signal LUT_gen20_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen20_block7_data : std_logic_vector(63 downto 0) := "1111000000001111111100000000111100001111111100000000111111110000";
   signal LUT_gen20_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen20_block8_data : std_logic_vector(63 downto 0) := "0101101010100101101001010101101001011010101001011010010101011010";
   signal LUT_gen20_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen20_block9_data : std_logic_vector(63 downto 0) := "1001100110011001100110011001100101100110011001100110011001100110";
   signal LUT_gen20_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen20_block10_data : std_logic_vector(63 downto 0) := "0000111100001111111100001111000000001111000011111111000011110000";
   signal LUT_gen20_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen20_block11_data : std_logic_vector(63 downto 0) := "1100001100111100001111001100001100111100110000111100001100111100";
   signal LUT_gen20_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen20_block12_data : std_logic_vector(63 downto 0) := "1111111100000000111111110000000011111111000000001111111100000000";
   signal LUT_gen20_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen20_block13_data : std_logic_vector(63 downto 0) := "1001011001101001100101100110100101101001100101100110100110010110";
   signal LUT_gen20_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen20_block14_data : std_logic_vector(63 downto 0) := "1111000011110000111100001111000011110000111100001111000011110000";
   signal LUT_gen20_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen20_block15_data : std_logic_vector(63 downto 0) := "0011110000111100110000111100001111000011110000110011110000111100";
   signal LUT_gen21 : std_logic_vector(15 downto 0);
   signal LUT_gen21_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen21_block0_data : std_logic_vector(63 downto 0) := "1001100101100110011001101001100101100110100110011001100101100110";
   signal LUT_gen21_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen21_block1_data : std_logic_vector(63 downto 0) := "1100001111000011110000111100001100111100001111000011110000111100";
   signal LUT_gen21_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen21_block2_data : std_logic_vector(63 downto 0) := "1100110011001100110011001100110011001100110011001100110011001100";
   signal LUT_gen21_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen21_block3_data : std_logic_vector(63 downto 0) := "0000000011111111000000001111111111111111000000001111111100000000";
   signal LUT_gen21_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen21_block4_data : std_logic_vector(63 downto 0) := "1010101001010101010101011010101010101010010101010101010110101010";
   signal LUT_gen21_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen21_block5_data : std_logic_vector(63 downto 0) := "1001011001101001100101100110100101101001100101100110100110010110";
   signal LUT_gen21_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen21_block6_data : std_logic_vector(63 downto 0) := "0110011010011001100110010110011001100110100110011001100101100110";
   signal LUT_gen21_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen21_block7_data : std_logic_vector(63 downto 0) := "0011001111001100001100111100110000110011110011000011001111001100";
   signal LUT_gen21_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen21_block8_data : std_logic_vector(63 downto 0) := "1111111111111111111111111111111100000000000000000000000000000000";
   signal LUT_gen21_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen21_block9_data : std_logic_vector(63 downto 0) := "1100001111000011110000111100001100111100001111000011110000111100";
   signal LUT_gen21_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen21_block10_data : std_logic_vector(63 downto 0) := "0101101010100101101001010101101001011010101001011010010101011010";
   signal LUT_gen21_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen21_block11_data : std_logic_vector(63 downto 0) := "1001100101100110100110010110011010011001011001101001100101100110";
   signal LUT_gen21_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen21_block12_data : std_logic_vector(63 downto 0) := "1111111111111111000000000000000011111111111111110000000000000000";
   signal LUT_gen21_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen21_block13_data : std_logic_vector(63 downto 0) := "1100110000110011001100111100110011001100001100110011001111001100";
   signal LUT_gen21_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen21_block14_data : std_logic_vector(63 downto 0) := "1111000011110000111100001111000011110000111100001111000011110000";
   signal LUT_gen21_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen21_block15_data : std_logic_vector(63 downto 0) := "0101101010100101010110101010010110100101010110101010010101011010";
   signal LUT_gen22 : std_logic_vector(15 downto 0);
   signal LUT_gen22_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen22_block0_data : std_logic_vector(63 downto 0) := "1111000000001111111100000000111100001111111100000000111111110000";
   signal LUT_gen22_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen22_block1_data : std_logic_vector(63 downto 0) := "1111000011110000000011110000111100001111000011111111000011110000";
   signal LUT_gen22_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen22_block2_data : std_logic_vector(63 downto 0) := "1010101010101010010101010101010101010101010101011010101010101010";
   signal LUT_gen22_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen22_block3_data : std_logic_vector(63 downto 0) := "1100001111000011001111000011110011000011110000110011110000111100";
   signal LUT_gen22_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen22_block4_data : std_logic_vector(63 downto 0) := "1001100101100110011001101001100101100110100110011001100101100110";
   signal LUT_gen22_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen22_block5_data : std_logic_vector(63 downto 0) := "0110011001100110100110011001100110011001100110010110011001100110";
   signal LUT_gen22_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen22_block6_data : std_logic_vector(63 downto 0) := "0011001100110011110011001100110000110011001100111100110011001100";
   signal LUT_gen22_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen22_block7_data : std_logic_vector(63 downto 0) := "1001011010010110100101101001011010010110100101101001011010010110";
   signal LUT_gen22_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen22_block8_data : std_logic_vector(63 downto 0) := "0110011010011001100110010110011001100110100110011001100101100110";
   signal LUT_gen22_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen22_block9_data : std_logic_vector(63 downto 0) := "0101101010100101010110101010010110100101010110101010010101011010";
   signal LUT_gen22_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen22_block10_data : std_logic_vector(63 downto 0) := "0110100110010110011010011001011001101001100101100110100110010110";
   signal LUT_gen22_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen22_block11_data : std_logic_vector(63 downto 0) := "0101010101010101010101010101010110101010101010101010101010101010";
   signal LUT_gen22_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen22_block12_data : std_logic_vector(63 downto 0) := "0101010101010101010101010101010110101010101010101010101010101010";
   signal LUT_gen22_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen22_block13_data : std_logic_vector(63 downto 0) := "0000000000000000111111111111111111111111111111110000000000000000";
   signal LUT_gen22_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen22_block14_data : std_logic_vector(63 downto 0) := "0101101001011010010110100101101001011010010110100101101001011010";
   signal LUT_gen22_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen22_block15_data : std_logic_vector(63 downto 0) := "0110011010011001100110010110011001100110100110011001100101100110";
   signal LUT_gen23 : std_logic_vector(15 downto 0);
   signal LUT_gen23_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen23_block0_data : std_logic_vector(63 downto 0) := "1010101001010101010101011010101010101010010101010101010110101010";
   signal LUT_gen23_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen23_block1_data : std_logic_vector(63 downto 0) := "1010101001010101101010100101010101010101101010100101010110101010";
   signal LUT_gen23_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen23_block2_data : std_logic_vector(63 downto 0) := "1001100110011001100110011001100101100110011001100110011001100110";
   signal LUT_gen23_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen23_block3_data : std_logic_vector(63 downto 0) := "0101101010100101010110101010010110100101010110101010010101011010";
   signal LUT_gen23_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen23_block4_data : std_logic_vector(63 downto 0) := "0011110000111100110000111100001111000011110000110011110000111100";
   signal LUT_gen23_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen23_block5_data : std_logic_vector(63 downto 0) := "0110100101101001011010010110100110010110100101101001011010010110";
   signal LUT_gen23_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen23_block6_data : std_logic_vector(63 downto 0) := "1010010110100101101001011010010101011010010110100101101001011010";
   signal LUT_gen23_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen23_block7_data : std_logic_vector(63 downto 0) := "1100001100111100110000110011110011000011001111001100001100111100";
   signal LUT_gen23_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen23_block8_data : std_logic_vector(63 downto 0) := "0011110000111100110000111100001111000011110000110011110000111100";
   signal LUT_gen23_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen23_block9_data : std_logic_vector(63 downto 0) := "1100110000110011001100111100110011001100001100110011001111001100";
   signal LUT_gen23_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen23_block10_data : std_logic_vector(63 downto 0) := "1001011001101001011010011001011010010110011010010110100110010110";
   signal LUT_gen23_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen23_block11_data : std_logic_vector(63 downto 0) := "1100110011001100110011001100110011001100110011001100110011001100";
   signal LUT_gen23_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen23_block12_data : std_logic_vector(63 downto 0) := "0110011001100110011001100110011001100110011001100110011001100110";
   signal LUT_gen23_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen23_block13_data : std_logic_vector(63 downto 0) := "0101010101010101010101010101010110101010101010101010101010101010";
   signal LUT_gen23_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen23_block14_data : std_logic_vector(63 downto 0) := "1001100101100110100110010110011010011001011001101001100101100110";
   signal LUT_gen23_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen23_block15_data : std_logic_vector(63 downto 0) := "0011110000111100110000111100001111000011110000110011110000111100";
   signal LUT_gen24 : std_logic_vector(15 downto 0);
   signal LUT_gen24_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen24_block0_data : std_logic_vector(63 downto 0) := "0000000011111111000000001111111111111111000000001111111100000000";
   signal LUT_gen24_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen24_block1_data : std_logic_vector(63 downto 0) := "0110011010011001011001101001100110011001011001101001100101100110";
   signal LUT_gen24_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen24_block2_data : std_logic_vector(63 downto 0) := "0110011001100110100110011001100110011001100110010110011001100110";
   signal LUT_gen24_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen24_block3_data : std_logic_vector(63 downto 0) := "0101101010100101101001010101101001011010101001011010010101011010";
   signal LUT_gen24_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen24_block4_data : std_logic_vector(63 downto 0) := "1010010110100101101001011010010101011010010110100101101001011010";
   signal LUT_gen24_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen24_block5_data : std_logic_vector(63 downto 0) := "0011001100110011001100110011001111001100110011001100110011001100";
   signal LUT_gen24_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen24_block6_data : std_logic_vector(63 downto 0) := "0011110011000011001111001100001111000011001111001100001100111100";
   signal LUT_gen24_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen24_block7_data : std_logic_vector(63 downto 0) := "1100001100111100110000110011110011000011001111001100001100111100";
   signal LUT_gen24_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen24_block8_data : std_logic_vector(63 downto 0) := "1001011010010110011010010110100101101001011010011001011010010110";
   signal LUT_gen24_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen24_block9_data : std_logic_vector(63 downto 0) := "1010010110100101010110100101101010100101101001010101101001011010";
   signal LUT_gen24_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen24_block10_data : std_logic_vector(63 downto 0) := "0011001111001100001100111100110000110011110011000011001111001100";
   signal LUT_gen24_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen24_block11_data : std_logic_vector(63 downto 0) := "0110011001100110100110011001100110011001100110010110011001100110";
   signal LUT_gen24_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen24_block12_data : std_logic_vector(63 downto 0) := "1001011010010110100101101001011010010110100101101001011010010110";
   signal LUT_gen24_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen24_block13_data : std_logic_vector(63 downto 0) := "0011110000111100001111000011110000111100001111000011110000111100";
   signal LUT_gen24_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen24_block14_data : std_logic_vector(63 downto 0) := "1100110000110011001100111100110011001100001100110011001111001100";
   signal LUT_gen24_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen24_block15_data : std_logic_vector(63 downto 0) := "0101101010100101010110101010010110100101010110101010010101011010";
   signal LUT_gen25 : std_logic_vector(15 downto 0);
   signal LUT_gen25_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen25_block0_data : std_logic_vector(63 downto 0) := "0011001111001100001100111100110000110011110011000011001111001100";
   signal LUT_gen25_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen25_block1_data : std_logic_vector(63 downto 0) := "0011110011000011001111001100001111000011001111001100001100111100";
   signal LUT_gen25_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen25_block2_data : std_logic_vector(63 downto 0) := "1001100110011001011001100110011010011001100110010110011001100110";
   signal LUT_gen25_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen25_block3_data : std_logic_vector(63 downto 0) := "1010010101011010010110101010010101011010101001011010010101011010";
   signal LUT_gen25_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen25_block4_data : std_logic_vector(63 downto 0) := "1100110011001100110011001100110011001100110011001100110011001100";
   signal LUT_gen25_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen25_block5_data : std_logic_vector(63 downto 0) := "0000000011111111000000001111111111111111000000001111111100000000";
   signal LUT_gen25_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen25_block6_data : std_logic_vector(63 downto 0) := "1111111100000000000000001111111100000000111111111111111100000000";
   signal LUT_gen25_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen25_block7_data : std_logic_vector(63 downto 0) := "1100001100111100110000110011110011000011001111001100001100111100";
   signal LUT_gen25_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen25_block8_data : std_logic_vector(63 downto 0) := "0101101001011010101001011010010110100101101001010101101001011010";
   signal LUT_gen25_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen25_block9_data : std_logic_vector(63 downto 0) := "1001100101100110100110010110011010011001011001101001100101100110";
   signal LUT_gen25_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen25_block10_data : std_logic_vector(63 downto 0) := "1111111111111111111111111111111100000000000000000000000000000000";
   signal LUT_gen25_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen25_block11_data : std_logic_vector(63 downto 0) := "0101010101010101101010101010101001010101010101011010101010101010";
   signal LUT_gen25_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen25_block12_data : std_logic_vector(63 downto 0) := "1100001100111100110000110011110011000011001111001100001100111100";
   signal LUT_gen25_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen25_block13_data : std_logic_vector(63 downto 0) := "1111111100000000111111110000000011111111000000001111111100000000";
   signal LUT_gen25_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen25_block14_data : std_logic_vector(63 downto 0) := "0101010110101010101010100101010110101010010101010101010110101010";
   signal LUT_gen25_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen25_block15_data : std_logic_vector(63 downto 0) := "0110011010011001100110010110011001100110100110011001100101100110";
   signal LUT_gen26 : std_logic_vector(15 downto 0);
   signal LUT_gen26_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen26_block0_data : std_logic_vector(63 downto 0) := "1010010110100101010110100101101010100101101001010101101001011010";
   signal LUT_gen26_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen26_block1_data : std_logic_vector(63 downto 0) := "1111000000001111000011111111000011110000000011110000111111110000";
   signal LUT_gen26_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen26_block2_data : std_logic_vector(63 downto 0) := "0110100101101001011010010110100110010110100101101001011010010110";
   signal LUT_gen26_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen26_block3_data : std_logic_vector(63 downto 0) := "0011001111001100110011000011001111001100001100110011001111001100";
   signal LUT_gen26_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen26_block4_data : std_logic_vector(63 downto 0) := "0101101001011010010110100101101001011010010110100101101001011010";
   signal LUT_gen26_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen26_block5_data : std_logic_vector(63 downto 0) := "0000111100001111111100001111000000001111000011111111000011110000";
   signal LUT_gen26_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen26_block6_data : std_logic_vector(63 downto 0) := "1010101010101010010101010101010101010101010101011010101010101010";
   signal LUT_gen26_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen26_block7_data : std_logic_vector(63 downto 0) := "0101101010100101101001010101101001011010101001011010010101011010";
   signal LUT_gen26_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen26_block8_data : std_logic_vector(63 downto 0) := "1100110000110011110011000011001100110011110011000011001111001100";
   signal LUT_gen26_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen26_block9_data : std_logic_vector(63 downto 0) := "0110100101101001100101101001011001101001011010011001011010010110";
   signal LUT_gen26_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen26_block11_data : std_logic_vector(63 downto 0) := "1001100110011001100110011001100101100110011001100110011001100110";
   signal LUT_gen26_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen26_block12_data : std_logic_vector(63 downto 0) := "1111000000001111000011111111000011110000000011110000111111110000";
   signal LUT_gen26_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen26_block13_data : std_logic_vector(63 downto 0) := "1111111111111111000000000000000011111111111111110000000000000000";
   signal LUT_gen26_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen26_block14_data : std_logic_vector(63 downto 0) := "1100110011001100001100110011001100110011001100111100110011001100";
   signal LUT_gen26_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen26_block15_data : std_logic_vector(63 downto 0) := "1001011010010110011010010110100101101001011010011001011010010110";
   signal LUT_gen27 : std_logic_vector(15 downto 0);
   signal LUT_gen27_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen27_block0_data : std_logic_vector(63 downto 0) := "1010101010101010010101010101010101010101010101011010101010101010";
   signal LUT_gen27_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen27_block1_data : std_logic_vector(63 downto 0) := "1010101010101010101010101010101010101010101010101010101010101010";
   signal LUT_gen27_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen27_block2_data : std_logic_vector(63 downto 0) := "0011001111001100110011000011001111001100001100110011001111001100";
   signal LUT_gen27_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen27_block3_data : std_logic_vector(63 downto 0) := "0110011001100110100110011001100110011001100110010110011001100110";
   signal LUT_gen27_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen27_block4_data : std_logic_vector(63 downto 0) := "0110011001100110011001100110011001100110011001100110011001100110";
   signal LUT_gen27_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen27_block5_data : std_logic_vector(63 downto 0) := "0101101001011010010110100101101001011010010110100101101001011010";
   signal LUT_gen27_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen27_block6_data : std_logic_vector(63 downto 0) := "1001011010010110100101101001011010010110100101101001011010010110";
   signal LUT_gen27_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen27_block7_data : std_logic_vector(63 downto 0) := "0000000011111111000000001111111111111111000000001111111100000000";
   signal LUT_gen27_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen27_block8_data : std_logic_vector(63 downto 0) := "0110100110010110011010011001011001101001100101100110100110010110";
   signal LUT_gen27_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen27_block9_data : std_logic_vector(63 downto 0) := "0110100110010110011010011001011001101001100101100110100110010110";
   signal LUT_gen27_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen27_block10_data : std_logic_vector(63 downto 0) := "1111000011110000000011110000111100001111000011111111000011110000";
   signal LUT_gen27_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen27_block11_data : std_logic_vector(63 downto 0) := "1010101010101010010101010101010101010101010101011010101010101010";
   signal LUT_gen27_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen27_block12_data : std_logic_vector(63 downto 0) := "1111111100000000000000001111111100000000111111111111111100000000";
   signal LUT_gen27_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen27_block13_data : std_logic_vector(63 downto 0) := "0000111100001111000011110000111111110000111100001111000011110000";
   signal LUT_gen27_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen27_block14_data : std_logic_vector(63 downto 0) := "1010101001010101101010100101010101010101101010100101010110101010";
   signal LUT_gen27_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen27_block15_data : std_logic_vector(63 downto 0) := "0011110011000011001111001100001111000011001111001100001100111100";
   signal LUT_gen28 : std_logic_vector(15 downto 0);
   signal LUT_gen28_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen28_block0_data : std_logic_vector(63 downto 0) := "1111111100000000000000001111111100000000111111111111111100000000";
   signal LUT_gen28_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen28_block1_data : std_logic_vector(63 downto 0) := "0011001111001100110011000011001111001100001100110011001111001100";
   signal LUT_gen28_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen28_block3_data : std_logic_vector(63 downto 0) := "0101010101010101010101010101010110101010101010101010101010101010";
   signal LUT_gen28_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen28_block4_data : std_logic_vector(63 downto 0) := "0110100110010110011010011001011001101001100101100110100110010110";
   signal LUT_gen28_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen28_block5_data : std_logic_vector(63 downto 0) := "1001100110011001100110011001100101100110011001100110011001100110";
   signal LUT_gen28_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen28_block6_data : std_logic_vector(63 downto 0) := "0110011010011001011001101001100110011001011001101001100101100110";
   signal LUT_gen28_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen28_block7_data : std_logic_vector(63 downto 0) := "0110011001100110011001100110011001100110011001100110011001100110";
   signal LUT_gen28_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen28_block8_data : std_logic_vector(63 downto 0) := "1111000011110000111100001111000011110000111100001111000011110000";
   signal LUT_gen28_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen28_block9_data : std_logic_vector(63 downto 0) := "1100001100111100001111001100001100111100110000111100001100111100";
   signal LUT_gen28_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen28_block10_data : std_logic_vector(63 downto 0) := "1111000000001111000011111111000011110000000011110000111111110000";
   signal LUT_gen28_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen28_block11_data : std_logic_vector(63 downto 0) := "0000111100001111111100001111000000001111000011111111000011110000";
   signal LUT_gen28_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen28_block12_data : std_logic_vector(63 downto 0) := "0000000000000000111111111111111111111111111111110000000000000000";
   signal LUT_gen28_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen28_block13_data : std_logic_vector(63 downto 0) := "1010010101011010101001010101101010100101010110101010010101011010";
   signal LUT_gen28_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen28_block14_data : std_logic_vector(63 downto 0) := "0011110011000011110000110011110000111100110000111100001100111100";
   signal LUT_gen28_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen28_block15_data : std_logic_vector(63 downto 0) := "1111000000001111000011111111000011110000000011110000111111110000";
   signal LUT_gen29 : std_logic_vector(15 downto 0);
   signal LUT_gen29_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen29_block0_data : std_logic_vector(63 downto 0) := "0000000000000000111111111111111111111111111111110000000000000000";
   signal LUT_gen29_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen29_block1_data : std_logic_vector(63 downto 0) := "0101101001011010101001011010010110100101101001010101101001011010";
   signal LUT_gen29_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen29_block2_data : std_logic_vector(63 downto 0) := "1010101010101010101010101010101010101010101010101010101010101010";
   signal LUT_gen29_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen29_block3_data : std_logic_vector(63 downto 0) := "1100110011001100110011001100110011001100110011001100110011001100";
   signal LUT_gen29_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen29_block4_data : std_logic_vector(63 downto 0) := "1001011001101001011010011001011010010110011010010110100110010110";
   signal LUT_gen29_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen29_block5_data : std_logic_vector(63 downto 0) := "1100110011001100110011001100110011001100110011001100110011001100";
   signal LUT_gen29_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen29_block6_data : std_logic_vector(63 downto 0) := "0110100101101001100101101001011001101001011010011001011010010110";
   signal LUT_gen29_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen29_block7_data : std_logic_vector(63 downto 0) := "1001011010010110100101101001011010010110100101101001011010010110";
   signal LUT_gen29_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen29_block8_data : std_logic_vector(63 downto 0) := "1111111100000000111111110000000011111111000000001111111100000000";
   signal LUT_gen29_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen29_block9_data : std_logic_vector(63 downto 0) := "0000111111110000111100000000111111110000000011110000111111110000";
   signal LUT_gen29_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen29_block10_data : std_logic_vector(63 downto 0) := "0101010110101010101010100101010110101010010101010101010110101010";
   signal LUT_gen29_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen29_block11_data : std_logic_vector(63 downto 0) := "0000000011111111000000001111111111111111000000001111111100000000";
   signal LUT_gen29_block12_addr : std_logic_vector(5 downto 0);
   constant LUT_gen29_block12_data : std_logic_vector(63 downto 0) := "1111111111111111111111111111111100000000000000000000000000000000";
   signal LUT_gen29_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen29_block13_data : std_logic_vector(63 downto 0) := "0110011010011001100110010110011001100110100110011001100101100110";
   signal LUT_gen29_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen29_block14_data : std_logic_vector(63 downto 0) := "0000111111110000111100000000111111110000000011110000111111110000";
   signal LUT_gen29_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen29_block15_data : std_logic_vector(63 downto 0) := "1111111100000000000000001111111100000000111111111111111100000000";
   signal LUT_gen30 : std_logic_vector(15 downto 0);
   signal LUT_gen30_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen30_block0_data : std_logic_vector(63 downto 0) := "1001100101100110011001101001100101100110100110011001100101100110";
   signal LUT_gen30_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen30_block1_data : std_logic_vector(63 downto 0) := "0011001100110011110011001100110000110011001100111100110011001100";
   signal LUT_gen30_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen30_block2_data : std_logic_vector(63 downto 0) := "1001011010010110011010010110100101101001011010011001011010010110";
   signal LUT_gen30_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen30_block3_data : std_logic_vector(63 downto 0) := "1100110011001100110011001100110011001100110011001100110011001100";
   signal LUT_gen30_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen30_block4_data : std_logic_vector(63 downto 0) := "0011110000111100110000111100001111000011110000110011110000111100";
   signal LUT_gen30_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen30_block5_data : std_logic_vector(63 downto 0) := "0101101010100101010110101010010110100101010110101010010101011010";
   signal LUT_gen30_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen30_block6_data : std_logic_vector(63 downto 0) := "1001100101100110100110010110011010011001011001101001100101100110";
   signal LUT_gen30_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen30_block7_data : std_logic_vector(63 downto 0) := "0101101010100101101001010101101001011010101001011010010101011010";
   signal LUT_gen30_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen30_block8_data : std_logic_vector(63 downto 0) := "1001100101100110100110010110011010011001011001101001100101100110";
   signal LUT_gen30_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen30_block9_data : std_logic_vector(63 downto 0) := "0000000011111111111111110000000000000000111111111111111100000000";
   signal LUT_gen30_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen30_block10_data : std_logic_vector(63 downto 0) := "1001011010010110100101101001011010010110100101101001011010010110";
   signal LUT_gen30_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen30_block11_data : std_logic_vector(63 downto 0) := "1100001111000011110000111100001100111100001111000011110000111100";
   signal LUT_gen30_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen30_block13_data : std_logic_vector(63 downto 0) := "0110011001100110100110011001100110011001100110010110011001100110";
   signal LUT_gen30_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen30_block14_data : std_logic_vector(63 downto 0) := "0101101001011010101001011010010110100101101001010101101001011010";
   signal LUT_gen30_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen30_block15_data : std_logic_vector(63 downto 0) := "0000000000000000111111111111111111111111111111110000000000000000";
   signal LUT_gen31 : std_logic_vector(15 downto 0);
   signal LUT_gen31_block0_addr : std_logic_vector(5 downto 0);
   constant LUT_gen31_block0_data : std_logic_vector(63 downto 0) := "0101101010100101010110101010010110100101010110101010010101011010";
   signal LUT_gen31_block1_addr : std_logic_vector(5 downto 0);
   constant LUT_gen31_block1_data : std_logic_vector(63 downto 0) := "1111000000001111000011111111000011110000000011110000111111110000";
   signal LUT_gen31_block2_addr : std_logic_vector(5 downto 0);
   constant LUT_gen31_block2_data : std_logic_vector(63 downto 0) := "1100110000110011001100111100110011001100001100110011001111001100";
   signal LUT_gen31_block3_addr : std_logic_vector(5 downto 0);
   constant LUT_gen31_block3_data : std_logic_vector(63 downto 0) := "0110011001100110011001100110011001100110011001100110011001100110";
   signal LUT_gen31_block4_addr : std_logic_vector(5 downto 0);
   constant LUT_gen31_block4_data : std_logic_vector(63 downto 0) := "0000111100001111000011110000111111110000111100001111000011110000";
   signal LUT_gen31_block5_addr : std_logic_vector(5 downto 0);
   constant LUT_gen31_block5_data : std_logic_vector(63 downto 0) := "0011110000111100110000111100001111000011110000110011110000111100";
   signal LUT_gen31_block6_addr : std_logic_vector(5 downto 0);
   constant LUT_gen31_block6_data : std_logic_vector(63 downto 0) := "1100110011001100001100110011001100110011001100111100110011001100";
   signal LUT_gen31_block7_addr : std_logic_vector(5 downto 0);
   constant LUT_gen31_block7_data : std_logic_vector(63 downto 0) := "1010101001010101101010100101010101010101101010100101010110101010";
   signal LUT_gen31_block8_addr : std_logic_vector(5 downto 0);
   constant LUT_gen31_block8_data : std_logic_vector(63 downto 0) := "1010010101011010101001010101101010100101010110101010010101011010";
   signal LUT_gen31_block9_addr : std_logic_vector(5 downto 0);
   constant LUT_gen31_block9_data : std_logic_vector(63 downto 0) := "1111111111111111000000000000000011111111111111110000000000000000";
   signal LUT_gen31_block10_addr : std_logic_vector(5 downto 0);
   constant LUT_gen31_block10_data : std_logic_vector(63 downto 0) := "0011001111001100110011000011001111001100001100110011001111001100";
   signal LUT_gen31_block11_addr : std_logic_vector(5 downto 0);
   constant LUT_gen31_block11_data : std_logic_vector(63 downto 0) := "1001100101100110011001101001100101100110100110011001100101100110";
   signal LUT_gen31_block13_addr : std_logic_vector(5 downto 0);
   constant LUT_gen31_block13_data : std_logic_vector(63 downto 0) := "0011001100110011001100110011001111001100110011001100110011001100";
   signal LUT_gen31_block14_addr : std_logic_vector(5 downto 0);
   constant LUT_gen31_block14_data : std_logic_vector(63 downto 0) := "1100001111000011110000111100001100111100001111000011110000111100";
   signal LUT_gen31_block15_addr : std_logic_vector(5 downto 0);
   constant LUT_gen31_block15_data : std_logic_vector(63 downto 0) := "1111111111111111111111111111111100000000000000000000000000000000";

   signal valid_del1 : std_logic := '0';
begin
   
   process(clk)
   begin 
      if rising_edge(clk) then 
         valid_del1 <= valid_i;
         if valid_i = '1' then
            cur_state <= new_state;
         end if;
      end if;
   end process;
   
   state_o <= cur_state;
   new_state_o <= new_state;
   

   new_state(0) <= LUT_gen0(0) xor LUT_gen0(1) xor LUT_gen0(2) xor LUT_gen0(3) xor LUT_gen0(4) xor LUT_gen0(5) xor LUT_gen0(6) xor LUT_gen0(7) xor LUT_gen0(8) xor LUT_gen0(9) xor LUT_gen0(10) xor LUT_gen0(11) xor LUT_gen0(12) xor LUT_gen0(13) xor LUT_gen0(14) xor LUT_gen0(15);
   new_state(1) <= LUT_gen1(0) xor LUT_gen1(1) xor LUT_gen1(2) xor LUT_gen1(3) xor LUT_gen1(4) xor LUT_gen1(5) xor LUT_gen1(6) xor LUT_gen1(7) xor LUT_gen1(8) xor LUT_gen1(9) xor LUT_gen1(10) xor LUT_gen1(11) xor LUT_gen1(12) xor LUT_gen1(13) xor LUT_gen1(14) xor LUT_gen1(15);
   new_state(2) <= LUT_gen2(0) xor LUT_gen2(1) xor LUT_gen2(2) xor LUT_gen2(3) xor LUT_gen2(4) xor LUT_gen2(5) xor LUT_gen2(6) xor LUT_gen2(7) xor LUT_gen2(8) xor LUT_gen2(9) xor LUT_gen2(10) xor LUT_gen2(11) xor LUT_gen2(12) xor LUT_gen2(13) xor LUT_gen2(14) xor LUT_gen2(15);
   new_state(3) <= LUT_gen3(0) xor LUT_gen3(1) xor LUT_gen3(2) xor LUT_gen3(3) xor LUT_gen3(4) xor LUT_gen3(5) xor LUT_gen3(6) xor LUT_gen3(7) xor LUT_gen3(8) xor LUT_gen3(9) xor LUT_gen3(10) xor LUT_gen3(11) xor LUT_gen3(12) xor LUT_gen3(13) xor LUT_gen3(14) xor LUT_gen3(15);
   new_state(4) <= LUT_gen4(0) xor LUT_gen4(1) xor LUT_gen4(2) xor LUT_gen4(3) xor LUT_gen4(4) xor LUT_gen4(5) xor LUT_gen4(6) xor LUT_gen4(7) xor LUT_gen4(8) xor LUT_gen4(9) xor LUT_gen4(10) xor LUT_gen4(11) xor LUT_gen4(12) xor LUT_gen4(13) xor LUT_gen4(14) xor LUT_gen4(15);
   new_state(5) <= LUT_gen5(0) xor LUT_gen5(1) xor LUT_gen5(2) xor LUT_gen5(3) xor LUT_gen5(4) xor LUT_gen5(5) xor LUT_gen5(6) xor LUT_gen5(7) xor LUT_gen5(8) xor LUT_gen5(9) xor LUT_gen5(10) xor LUT_gen5(11) xor LUT_gen5(12) xor LUT_gen5(13) xor LUT_gen5(14) xor LUT_gen5(15);
   new_state(6) <= LUT_gen6(0) xor LUT_gen6(1) xor LUT_gen6(2) xor LUT_gen6(3) xor LUT_gen6(4) xor LUT_gen6(5) xor LUT_gen6(6) xor LUT_gen6(7) xor LUT_gen6(8) xor LUT_gen6(9) xor LUT_gen6(10) xor LUT_gen6(11) xor LUT_gen6(12) xor LUT_gen6(13) xor LUT_gen6(14) xor LUT_gen6(15);
   new_state(7) <= LUT_gen7(0) xor LUT_gen7(1) xor LUT_gen7(2) xor LUT_gen7(3) xor LUT_gen7(4) xor LUT_gen7(5) xor LUT_gen7(6) xor LUT_gen7(7) xor LUT_gen7(8) xor LUT_gen7(9) xor LUT_gen7(10) xor LUT_gen7(11) xor LUT_gen7(12) xor LUT_gen7(13) xor LUT_gen7(14) xor LUT_gen7(15);
   new_state(8) <= LUT_gen8(0) xor LUT_gen8(1) xor LUT_gen8(2) xor LUT_gen8(3) xor LUT_gen8(4) xor LUT_gen8(5) xor LUT_gen8(6) xor LUT_gen8(7) xor LUT_gen8(8) xor LUT_gen8(9) xor LUT_gen8(10) xor LUT_gen8(11) xor LUT_gen8(12) xor LUT_gen8(13) xor LUT_gen8(14) xor LUT_gen8(15);
   new_state(9) <= LUT_gen9(0) xor LUT_gen9(1) xor LUT_gen9(2) xor LUT_gen9(3) xor LUT_gen9(4) xor LUT_gen9(5) xor LUT_gen9(6) xor LUT_gen9(7) xor LUT_gen9(8) xor LUT_gen9(9) xor LUT_gen9(10) xor LUT_gen9(11) xor LUT_gen9(12) xor LUT_gen9(13) xor LUT_gen9(14) xor LUT_gen9(15);
   new_state(10) <= LUT_gen10(0) xor LUT_gen10(1) xor LUT_gen10(2) xor LUT_gen10(3) xor LUT_gen10(4) xor LUT_gen10(5) xor LUT_gen10(6) xor LUT_gen10(7) xor LUT_gen10(8) xor LUT_gen10(9) xor LUT_gen10(10) xor LUT_gen10(11) xor LUT_gen10(12) xor LUT_gen10(13) xor LUT_gen10(14) xor LUT_gen10(15);
   new_state(11) <= LUT_gen11(0) xor LUT_gen11(1) xor LUT_gen11(2) xor LUT_gen11(3) xor LUT_gen11(4) xor LUT_gen11(5) xor LUT_gen11(6) xor LUT_gen11(7) xor LUT_gen11(8) xor LUT_gen11(9) xor LUT_gen11(10) xor LUT_gen11(11) xor LUT_gen11(12) xor LUT_gen11(13) xor LUT_gen11(14) xor LUT_gen11(15);
   new_state(12) <= LUT_gen12(0) xor LUT_gen12(1) xor LUT_gen12(2) xor LUT_gen12(3) xor LUT_gen12(4) xor LUT_gen12(5) xor LUT_gen12(6) xor LUT_gen12(7) xor LUT_gen12(8) xor LUT_gen12(9) xor LUT_gen12(10) xor LUT_gen12(11) xor LUT_gen12(12) xor LUT_gen12(13) xor LUT_gen12(14) xor LUT_gen12(15);
   new_state(13) <= LUT_gen13(0) xor LUT_gen13(1) xor LUT_gen13(2) xor LUT_gen13(3) xor LUT_gen13(4) xor LUT_gen13(5) xor LUT_gen13(6) xor LUT_gen13(7) xor LUT_gen13(8) xor LUT_gen13(9) xor LUT_gen13(10) xor LUT_gen13(11) xor LUT_gen13(12) xor LUT_gen13(13) xor LUT_gen13(14) xor LUT_gen13(15);
   new_state(14) <= LUT_gen14(0) xor LUT_gen14(1) xor LUT_gen14(2) xor LUT_gen14(3) xor LUT_gen14(4) xor LUT_gen14(5) xor LUT_gen14(6) xor LUT_gen14(7) xor LUT_gen14(8) xor LUT_gen14(9) xor LUT_gen14(10) xor LUT_gen14(11) xor LUT_gen14(12) xor LUT_gen14(13) xor LUT_gen14(14) xor LUT_gen14(15);
   new_state(15) <= LUT_gen15(0) xor LUT_gen15(1) xor LUT_gen15(2) xor LUT_gen15(3) xor LUT_gen15(4) xor LUT_gen15(5) xor LUT_gen15(6) xor LUT_gen15(7) xor LUT_gen15(8) xor LUT_gen15(9) xor LUT_gen15(10) xor LUT_gen15(11) xor LUT_gen15(12) xor LUT_gen15(13) xor LUT_gen15(14) xor LUT_gen15(15);
   new_state(16) <= LUT_gen16(0) xor LUT_gen16(1) xor LUT_gen16(2) xor LUT_gen16(3) xor LUT_gen16(4) xor LUT_gen16(5) xor LUT_gen16(6) xor LUT_gen16(7) xor LUT_gen16(8) xor LUT_gen16(9) xor LUT_gen16(10) xor LUT_gen16(11) xor LUT_gen16(12) xor LUT_gen16(13) xor LUT_gen16(14) xor LUT_gen16(15);
   new_state(17) <= LUT_gen17(0) xor LUT_gen17(1) xor LUT_gen17(2) xor LUT_gen17(3) xor LUT_gen17(4) xor LUT_gen17(5) xor LUT_gen17(6) xor LUT_gen17(7) xor LUT_gen17(8) xor LUT_gen17(9) xor LUT_gen17(10) xor LUT_gen17(11) xor LUT_gen17(12) xor LUT_gen17(13) xor LUT_gen17(14) xor LUT_gen17(15);
   new_state(18) <= LUT_gen18(0) xor LUT_gen18(1) xor LUT_gen18(2) xor LUT_gen18(3) xor LUT_gen18(4) xor LUT_gen18(5) xor LUT_gen18(6) xor LUT_gen18(7) xor LUT_gen18(8) xor LUT_gen18(9) xor LUT_gen18(10) xor LUT_gen18(11) xor LUT_gen18(12) xor LUT_gen18(13) xor LUT_gen18(14) xor LUT_gen18(15);
   new_state(19) <= LUT_gen19(0) xor LUT_gen19(1) xor LUT_gen19(2) xor LUT_gen19(3) xor LUT_gen19(4) xor LUT_gen19(5) xor LUT_gen19(6) xor LUT_gen19(7) xor LUT_gen19(8) xor LUT_gen19(9) xor LUT_gen19(10) xor LUT_gen19(11) xor LUT_gen19(12) xor LUT_gen19(13) xor LUT_gen19(14) xor LUT_gen19(15);
   new_state(20) <= LUT_gen20(0) xor LUT_gen20(1) xor LUT_gen20(2) xor LUT_gen20(3) xor LUT_gen20(4) xor LUT_gen20(5) xor LUT_gen20(6) xor LUT_gen20(7) xor LUT_gen20(8) xor LUT_gen20(9) xor LUT_gen20(10) xor LUT_gen20(11) xor LUT_gen20(12) xor LUT_gen20(13) xor LUT_gen20(14) xor LUT_gen20(15);
   new_state(21) <= LUT_gen21(0) xor LUT_gen21(1) xor LUT_gen21(2) xor LUT_gen21(3) xor LUT_gen21(4) xor LUT_gen21(5) xor LUT_gen21(6) xor LUT_gen21(7) xor LUT_gen21(8) xor LUT_gen21(9) xor LUT_gen21(10) xor LUT_gen21(11) xor LUT_gen21(12) xor LUT_gen21(13) xor LUT_gen21(14) xor LUT_gen21(15);
   new_state(22) <= LUT_gen22(0) xor LUT_gen22(1) xor LUT_gen22(2) xor LUT_gen22(3) xor LUT_gen22(4) xor LUT_gen22(5) xor LUT_gen22(6) xor LUT_gen22(7) xor LUT_gen22(8) xor LUT_gen22(9) xor LUT_gen22(10) xor LUT_gen22(11) xor LUT_gen22(12) xor LUT_gen22(13) xor LUT_gen22(14) xor LUT_gen22(15);
   new_state(23) <= LUT_gen23(0) xor LUT_gen23(1) xor LUT_gen23(2) xor LUT_gen23(3) xor LUT_gen23(4) xor LUT_gen23(5) xor LUT_gen23(6) xor LUT_gen23(7) xor LUT_gen23(8) xor LUT_gen23(9) xor LUT_gen23(10) xor LUT_gen23(11) xor LUT_gen23(12) xor LUT_gen23(13) xor LUT_gen23(14) xor LUT_gen23(15);
   new_state(24) <= LUT_gen24(0) xor LUT_gen24(1) xor LUT_gen24(2) xor LUT_gen24(3) xor LUT_gen24(4) xor LUT_gen24(5) xor LUT_gen24(6) xor LUT_gen24(7) xor LUT_gen24(8) xor LUT_gen24(9) xor LUT_gen24(10) xor LUT_gen24(11) xor LUT_gen24(12) xor LUT_gen24(13) xor LUT_gen24(14) xor LUT_gen24(15);
   new_state(25) <= LUT_gen25(0) xor LUT_gen25(1) xor LUT_gen25(2) xor LUT_gen25(3) xor LUT_gen25(4) xor LUT_gen25(5) xor LUT_gen25(6) xor LUT_gen25(7) xor LUT_gen25(8) xor LUT_gen25(9) xor LUT_gen25(10) xor LUT_gen25(11) xor LUT_gen25(12) xor LUT_gen25(13) xor LUT_gen25(14) xor LUT_gen25(15);
   new_state(26) <= LUT_gen26(0) xor LUT_gen26(1) xor LUT_gen26(2) xor LUT_gen26(3) xor LUT_gen26(4) xor LUT_gen26(5) xor LUT_gen26(6) xor LUT_gen26(7) xor LUT_gen26(8) xor LUT_gen26(9) xor LUT_gen26(10) xor LUT_gen26(11) xor LUT_gen26(12) xor LUT_gen26(13) xor LUT_gen26(14) xor LUT_gen26(15);
   new_state(27) <= LUT_gen27(0) xor LUT_gen27(1) xor LUT_gen27(2) xor LUT_gen27(3) xor LUT_gen27(4) xor LUT_gen27(5) xor LUT_gen27(6) xor LUT_gen27(7) xor LUT_gen27(8) xor LUT_gen27(9) xor LUT_gen27(10) xor LUT_gen27(11) xor LUT_gen27(12) xor LUT_gen27(13) xor LUT_gen27(14) xor LUT_gen27(15);
   new_state(28) <= LUT_gen28(0) xor LUT_gen28(1) xor LUT_gen28(2) xor LUT_gen28(3) xor LUT_gen28(4) xor LUT_gen28(5) xor LUT_gen28(6) xor LUT_gen28(7) xor LUT_gen28(8) xor LUT_gen28(9) xor LUT_gen28(10) xor LUT_gen28(11) xor LUT_gen28(12) xor LUT_gen28(13) xor LUT_gen28(14) xor LUT_gen28(15);
   new_state(29) <= LUT_gen29(0) xor LUT_gen29(1) xor LUT_gen29(2) xor LUT_gen29(3) xor LUT_gen29(4) xor LUT_gen29(5) xor LUT_gen29(6) xor LUT_gen29(7) xor LUT_gen29(8) xor LUT_gen29(9) xor LUT_gen29(10) xor LUT_gen29(11) xor LUT_gen29(12) xor LUT_gen29(13) xor LUT_gen29(14) xor LUT_gen29(15);
   new_state(30) <= LUT_gen30(0) xor LUT_gen30(1) xor LUT_gen30(2) xor LUT_gen30(3) xor LUT_gen30(4) xor LUT_gen30(5) xor LUT_gen30(6) xor LUT_gen30(7) xor LUT_gen30(8) xor LUT_gen30(9) xor LUT_gen30(10) xor LUT_gen30(11) xor LUT_gen30(12) xor LUT_gen30(13) xor LUT_gen30(14) xor LUT_gen30(15);
   new_state(31) <= LUT_gen31(0) xor LUT_gen31(1) xor LUT_gen31(2) xor LUT_gen31(3) xor LUT_gen31(4) xor LUT_gen31(5) xor LUT_gen31(6) xor LUT_gen31(7) xor LUT_gen31(8) xor LUT_gen31(9) xor LUT_gen31(10) xor LUT_gen31(11) xor LUT_gen31(12) xor LUT_gen31(13) xor LUT_gen31(14) xor LUT_gen31(15);


   allbits <= data_i & cur_state when sof_i = '0' else data_i & x"ffffffff"; -- Concatenate the data bits and state bits to make selecting them easier 
   LUT_gen0_block0_addr <= allbits(5 downto 0);
   LUT_gen0(0) <= LUT_gen0_block0_data(to_integer(unsigned(LUT_gen0_block0_addr)));
   LUT_gen0_block1_addr <= allbits(11 downto 6);
   LUT_gen0(1) <= LUT_gen0_block1_data(to_integer(unsigned(LUT_gen0_block1_addr)));
   LUT_gen0_block2_addr <= allbits(17 downto 12);
   LUT_gen0(2) <= LUT_gen0_block2_data(to_integer(unsigned(LUT_gen0_block2_addr)));
   LUT_gen0_block3_addr <= allbits(23 downto 18);
   LUT_gen0(3) <= LUT_gen0_block3_data(to_integer(unsigned(LUT_gen0_block3_addr)));
   LUT_gen0_block4_addr <= allbits(29 downto 24);
   LUT_gen0(4) <= LUT_gen0_block4_data(to_integer(unsigned(LUT_gen0_block4_addr)));
   LUT_gen0_block5_addr <= allbits(35 downto 30);
   LUT_gen0(5) <= LUT_gen0_block5_data(to_integer(unsigned(LUT_gen0_block5_addr)));
   LUT_gen0_block6_addr <= allbits(41 downto 36);
   LUT_gen0(6) <= LUT_gen0_block6_data(to_integer(unsigned(LUT_gen0_block6_addr)));
   LUT_gen0_block7_addr <= allbits(47 downto 42);
   LUT_gen0(7) <= LUT_gen0_block7_data(to_integer(unsigned(LUT_gen0_block7_addr)));
   LUT_gen0_block8_addr <= allbits(53 downto 48);
   LUT_gen0(8) <= LUT_gen0_block8_data(to_integer(unsigned(LUT_gen0_block8_addr)));
   LUT_gen0_block9_addr <= allbits(59 downto 54);
   LUT_gen0(9) <= LUT_gen0_block9_data(to_integer(unsigned(LUT_gen0_block9_addr)));
   LUT_gen0_block10_addr <= allbits(65 downto 60);
   LUT_gen0(10) <= LUT_gen0_block10_data(to_integer(unsigned(LUT_gen0_block10_addr)));
   LUT_gen0_block11_addr <= allbits(71 downto 66);
   LUT_gen0(11) <= LUT_gen0_block11_data(to_integer(unsigned(LUT_gen0_block11_addr)));
   LUT_gen0_block12_addr <= allbits(77 downto 72);
   LUT_gen0(12) <= LUT_gen0_block12_data(to_integer(unsigned(LUT_gen0_block12_addr)));
   LUT_gen0_block13_addr <= allbits(83 downto 78);
   LUT_gen0(13) <= LUT_gen0_block13_data(to_integer(unsigned(LUT_gen0_block13_addr)));
   LUT_gen0_block14_addr <= allbits(89 downto 84);
   LUT_gen0(14) <= LUT_gen0_block14_data(to_integer(unsigned(LUT_gen0_block14_addr)));
   LUT_gen0_block15_addr <= allbits(95 downto 90);
   LUT_gen0(15) <= LUT_gen0_block15_data(to_integer(unsigned(LUT_gen0_block15_addr)));
   LUT_gen1_block0_addr <= allbits(5 downto 0);
   LUT_gen1(0) <= LUT_gen1_block0_data(to_integer(unsigned(LUT_gen1_block0_addr)));
   LUT_gen1_block1_addr <= allbits(11 downto 6);
   LUT_gen1(1) <= LUT_gen1_block1_data(to_integer(unsigned(LUT_gen1_block1_addr)));
   LUT_gen1_block2_addr <= allbits(17 downto 12);
   LUT_gen1(2) <= LUT_gen1_block2_data(to_integer(unsigned(LUT_gen1_block2_addr)));
   LUT_gen1_block3_addr <= allbits(23 downto 18);
   LUT_gen1(3) <= LUT_gen1_block3_data(to_integer(unsigned(LUT_gen1_block3_addr)));
   LUT_gen1_block4_addr <= allbits(29 downto 24);
   LUT_gen1(4) <= LUT_gen1_block4_data(to_integer(unsigned(LUT_gen1_block4_addr)));
   LUT_gen1_block5_addr <= allbits(35 downto 30);
   LUT_gen1(5) <= LUT_gen1_block5_data(to_integer(unsigned(LUT_gen1_block5_addr)));
   LUT_gen1_block6_addr <= allbits(41 downto 36);
   LUT_gen1(6) <= LUT_gen1_block6_data(to_integer(unsigned(LUT_gen1_block6_addr)));
   LUT_gen1_block7_addr <= allbits(47 downto 42);
   LUT_gen1(7) <= LUT_gen1_block7_data(to_integer(unsigned(LUT_gen1_block7_addr)));
   LUT_gen1_block8_addr <= allbits(53 downto 48);
   LUT_gen1(8) <= LUT_gen1_block8_data(to_integer(unsigned(LUT_gen1_block8_addr)));
   LUT_gen1(9) <= '0';
   LUT_gen1_block10_addr <= allbits(65 downto 60);
   LUT_gen1(10) <= LUT_gen1_block10_data(to_integer(unsigned(LUT_gen1_block10_addr)));
   LUT_gen1_block11_addr <= allbits(71 downto 66);
   LUT_gen1(11) <= LUT_gen1_block11_data(to_integer(unsigned(LUT_gen1_block11_addr)));
   LUT_gen1_block12_addr <= allbits(77 downto 72);
   LUT_gen1(12) <= LUT_gen1_block12_data(to_integer(unsigned(LUT_gen1_block12_addr)));
   LUT_gen1_block13_addr <= allbits(83 downto 78);
   LUT_gen1(13) <= LUT_gen1_block13_data(to_integer(unsigned(LUT_gen1_block13_addr)));
   LUT_gen1_block14_addr <= allbits(89 downto 84);
   LUT_gen1(14) <= LUT_gen1_block14_data(to_integer(unsigned(LUT_gen1_block14_addr)));
   LUT_gen1_block15_addr <= allbits(95 downto 90);
   LUT_gen1(15) <= LUT_gen1_block15_data(to_integer(unsigned(LUT_gen1_block15_addr)));
   LUT_gen2_block0_addr <= allbits(5 downto 0);
   LUT_gen2(0) <= LUT_gen2_block0_data(to_integer(unsigned(LUT_gen2_block0_addr)));
   LUT_gen2_block1_addr <= allbits(11 downto 6);
   LUT_gen2(1) <= LUT_gen2_block1_data(to_integer(unsigned(LUT_gen2_block1_addr)));
   LUT_gen2_block2_addr <= allbits(17 downto 12);
   LUT_gen2(2) <= LUT_gen2_block2_data(to_integer(unsigned(LUT_gen2_block2_addr)));
   LUT_gen2_block3_addr <= allbits(23 downto 18);
   LUT_gen2(3) <= LUT_gen2_block3_data(to_integer(unsigned(LUT_gen2_block3_addr)));
   LUT_gen2_block4_addr <= allbits(29 downto 24);
   LUT_gen2(4) <= LUT_gen2_block4_data(to_integer(unsigned(LUT_gen2_block4_addr)));
   LUT_gen2_block5_addr <= allbits(35 downto 30);
   LUT_gen2(5) <= LUT_gen2_block5_data(to_integer(unsigned(LUT_gen2_block5_addr)));
   LUT_gen2_block6_addr <= allbits(41 downto 36);
   LUT_gen2(6) <= LUT_gen2_block6_data(to_integer(unsigned(LUT_gen2_block6_addr)));
   LUT_gen2_block7_addr <= allbits(47 downto 42);
   LUT_gen2(7) <= LUT_gen2_block7_data(to_integer(unsigned(LUT_gen2_block7_addr)));
   LUT_gen2_block8_addr <= allbits(53 downto 48);
   LUT_gen2(8) <= LUT_gen2_block8_data(to_integer(unsigned(LUT_gen2_block8_addr)));
   LUT_gen2_block9_addr <= allbits(59 downto 54);
   LUT_gen2(9) <= LUT_gen2_block9_data(to_integer(unsigned(LUT_gen2_block9_addr)));
   LUT_gen2_block10_addr <= allbits(65 downto 60);
   LUT_gen2(10) <= LUT_gen2_block10_data(to_integer(unsigned(LUT_gen2_block10_addr)));
   LUT_gen2_block11_addr <= allbits(71 downto 66);
   LUT_gen2(11) <= LUT_gen2_block11_data(to_integer(unsigned(LUT_gen2_block11_addr)));
   LUT_gen2_block12_addr <= allbits(77 downto 72);
   LUT_gen2(12) <= LUT_gen2_block12_data(to_integer(unsigned(LUT_gen2_block12_addr)));
   LUT_gen2_block13_addr <= allbits(83 downto 78);
   LUT_gen2(13) <= LUT_gen2_block13_data(to_integer(unsigned(LUT_gen2_block13_addr)));
   LUT_gen2_block14_addr <= allbits(89 downto 84);
   LUT_gen2(14) <= LUT_gen2_block14_data(to_integer(unsigned(LUT_gen2_block14_addr)));
   LUT_gen2_block15_addr <= allbits(95 downto 90);
   LUT_gen2(15) <= LUT_gen2_block15_data(to_integer(unsigned(LUT_gen2_block15_addr)));
   LUT_gen3_block0_addr <= allbits(5 downto 0);
   LUT_gen3(0) <= LUT_gen3_block0_data(to_integer(unsigned(LUT_gen3_block0_addr)));
   LUT_gen3_block1_addr <= allbits(11 downto 6);
   LUT_gen3(1) <= LUT_gen3_block1_data(to_integer(unsigned(LUT_gen3_block1_addr)));
   LUT_gen3_block2_addr <= allbits(17 downto 12);
   LUT_gen3(2) <= LUT_gen3_block2_data(to_integer(unsigned(LUT_gen3_block2_addr)));
   LUT_gen3_block3_addr <= allbits(23 downto 18);
   LUT_gen3(3) <= LUT_gen3_block3_data(to_integer(unsigned(LUT_gen3_block3_addr)));
   LUT_gen3(4) <= '0';
   LUT_gen3_block5_addr <= allbits(35 downto 30);
   LUT_gen3(5) <= LUT_gen3_block5_data(to_integer(unsigned(LUT_gen3_block5_addr)));
   LUT_gen3_block6_addr <= allbits(41 downto 36);
   LUT_gen3(6) <= LUT_gen3_block6_data(to_integer(unsigned(LUT_gen3_block6_addr)));
   LUT_gen3_block7_addr <= allbits(47 downto 42);
   LUT_gen3(7) <= LUT_gen3_block7_data(to_integer(unsigned(LUT_gen3_block7_addr)));
   LUT_gen3_block8_addr <= allbits(53 downto 48);
   LUT_gen3(8) <= LUT_gen3_block8_data(to_integer(unsigned(LUT_gen3_block8_addr)));
   LUT_gen3_block9_addr <= allbits(59 downto 54);
   LUT_gen3(9) <= LUT_gen3_block9_data(to_integer(unsigned(LUT_gen3_block9_addr)));
   LUT_gen3_block10_addr <= allbits(65 downto 60);
   LUT_gen3(10) <= LUT_gen3_block10_data(to_integer(unsigned(LUT_gen3_block10_addr)));
   LUT_gen3_block11_addr <= allbits(71 downto 66);
   LUT_gen3(11) <= LUT_gen3_block11_data(to_integer(unsigned(LUT_gen3_block11_addr)));
   LUT_gen3_block12_addr <= allbits(77 downto 72);
   LUT_gen3(12) <= LUT_gen3_block12_data(to_integer(unsigned(LUT_gen3_block12_addr)));
   LUT_gen3_block13_addr <= allbits(83 downto 78);
   LUT_gen3(13) <= LUT_gen3_block13_data(to_integer(unsigned(LUT_gen3_block13_addr)));
   LUT_gen3_block14_addr <= allbits(89 downto 84);
   LUT_gen3(14) <= LUT_gen3_block14_data(to_integer(unsigned(LUT_gen3_block14_addr)));
   LUT_gen3_block15_addr <= allbits(95 downto 90);
   LUT_gen3(15) <= LUT_gen3_block15_data(to_integer(unsigned(LUT_gen3_block15_addr)));
   LUT_gen4_block0_addr <= allbits(5 downto 0);
   LUT_gen4(0) <= LUT_gen4_block0_data(to_integer(unsigned(LUT_gen4_block0_addr)));
   LUT_gen4_block1_addr <= allbits(11 downto 6);
   LUT_gen4(1) <= LUT_gen4_block1_data(to_integer(unsigned(LUT_gen4_block1_addr)));
   LUT_gen4_block2_addr <= allbits(17 downto 12);
   LUT_gen4(2) <= LUT_gen4_block2_data(to_integer(unsigned(LUT_gen4_block2_addr)));
   LUT_gen4_block3_addr <= allbits(23 downto 18);
   LUT_gen4(3) <= LUT_gen4_block3_data(to_integer(unsigned(LUT_gen4_block3_addr)));
   LUT_gen4_block4_addr <= allbits(29 downto 24);
   LUT_gen4(4) <= LUT_gen4_block4_data(to_integer(unsigned(LUT_gen4_block4_addr)));
   LUT_gen4_block5_addr <= allbits(35 downto 30);
   LUT_gen4(5) <= LUT_gen4_block5_data(to_integer(unsigned(LUT_gen4_block5_addr)));
   LUT_gen4_block6_addr <= allbits(41 downto 36);
   LUT_gen4(6) <= LUT_gen4_block6_data(to_integer(unsigned(LUT_gen4_block6_addr)));
   LUT_gen4_block7_addr <= allbits(47 downto 42);
   LUT_gen4(7) <= LUT_gen4_block7_data(to_integer(unsigned(LUT_gen4_block7_addr)));
   LUT_gen4_block8_addr <= allbits(53 downto 48);
   LUT_gen4(8) <= LUT_gen4_block8_data(to_integer(unsigned(LUT_gen4_block8_addr)));
   LUT_gen4_block9_addr <= allbits(59 downto 54);
   LUT_gen4(9) <= LUT_gen4_block9_data(to_integer(unsigned(LUT_gen4_block9_addr)));
   LUT_gen4_block10_addr <= allbits(65 downto 60);
   LUT_gen4(10) <= LUT_gen4_block10_data(to_integer(unsigned(LUT_gen4_block10_addr)));
   LUT_gen4_block11_addr <= allbits(71 downto 66);
   LUT_gen4(11) <= LUT_gen4_block11_data(to_integer(unsigned(LUT_gen4_block11_addr)));
   LUT_gen4_block12_addr <= allbits(77 downto 72);
   LUT_gen4(12) <= LUT_gen4_block12_data(to_integer(unsigned(LUT_gen4_block12_addr)));
   LUT_gen4(13) <= '0';
   LUT_gen4_block14_addr <= allbits(89 downto 84);
   LUT_gen4(14) <= LUT_gen4_block14_data(to_integer(unsigned(LUT_gen4_block14_addr)));
   LUT_gen4_block15_addr <= allbits(95 downto 90);
   LUT_gen4(15) <= LUT_gen4_block15_data(to_integer(unsigned(LUT_gen4_block15_addr)));
   LUT_gen5_block0_addr <= allbits(5 downto 0);
   LUT_gen5(0) <= LUT_gen5_block0_data(to_integer(unsigned(LUT_gen5_block0_addr)));
   LUT_gen5_block1_addr <= allbits(11 downto 6);
   LUT_gen5(1) <= LUT_gen5_block1_data(to_integer(unsigned(LUT_gen5_block1_addr)));
   LUT_gen5_block2_addr <= allbits(17 downto 12);
   LUT_gen5(2) <= LUT_gen5_block2_data(to_integer(unsigned(LUT_gen5_block2_addr)));
   LUT_gen5_block3_addr <= allbits(23 downto 18);
   LUT_gen5(3) <= LUT_gen5_block3_data(to_integer(unsigned(LUT_gen5_block3_addr)));
   LUT_gen5_block4_addr <= allbits(29 downto 24);
   LUT_gen5(4) <= LUT_gen5_block4_data(to_integer(unsigned(LUT_gen5_block4_addr)));
   LUT_gen5_block5_addr <= allbits(35 downto 30);
   LUT_gen5(5) <= LUT_gen5_block5_data(to_integer(unsigned(LUT_gen5_block5_addr)));
   LUT_gen5_block6_addr <= allbits(41 downto 36);
   LUT_gen5(6) <= LUT_gen5_block6_data(to_integer(unsigned(LUT_gen5_block6_addr)));
   LUT_gen5_block7_addr <= allbits(47 downto 42);
   LUT_gen5(7) <= LUT_gen5_block7_data(to_integer(unsigned(LUT_gen5_block7_addr)));
   LUT_gen5_block8_addr <= allbits(53 downto 48);
   LUT_gen5(8) <= LUT_gen5_block8_data(to_integer(unsigned(LUT_gen5_block8_addr)));
   LUT_gen5_block9_addr <= allbits(59 downto 54);
   LUT_gen5(9) <= LUT_gen5_block9_data(to_integer(unsigned(LUT_gen5_block9_addr)));
   LUT_gen5_block10_addr <= allbits(65 downto 60);
   LUT_gen5(10) <= LUT_gen5_block10_data(to_integer(unsigned(LUT_gen5_block10_addr)));
   LUT_gen5_block11_addr <= allbits(71 downto 66);
   LUT_gen5(11) <= LUT_gen5_block11_data(to_integer(unsigned(LUT_gen5_block11_addr)));
   LUT_gen5_block12_addr <= allbits(77 downto 72);
   LUT_gen5(12) <= LUT_gen5_block12_data(to_integer(unsigned(LUT_gen5_block12_addr)));
   LUT_gen5(13) <= '0';
   LUT_gen5_block14_addr <= allbits(89 downto 84);
   LUT_gen5(14) <= LUT_gen5_block14_data(to_integer(unsigned(LUT_gen5_block14_addr)));
   LUT_gen5_block15_addr <= allbits(95 downto 90);
   LUT_gen5(15) <= LUT_gen5_block15_data(to_integer(unsigned(LUT_gen5_block15_addr)));
   LUT_gen6_block0_addr <= allbits(5 downto 0);
   LUT_gen6(0) <= LUT_gen6_block0_data(to_integer(unsigned(LUT_gen6_block0_addr)));
   LUT_gen6_block1_addr <= allbits(11 downto 6);
   LUT_gen6(1) <= LUT_gen6_block1_data(to_integer(unsigned(LUT_gen6_block1_addr)));
   LUT_gen6_block2_addr <= allbits(17 downto 12);
   LUT_gen6(2) <= LUT_gen6_block2_data(to_integer(unsigned(LUT_gen6_block2_addr)));
   LUT_gen6_block3_addr <= allbits(23 downto 18);
   LUT_gen6(3) <= LUT_gen6_block3_data(to_integer(unsigned(LUT_gen6_block3_addr)));
   LUT_gen6_block4_addr <= allbits(29 downto 24);
   LUT_gen6(4) <= LUT_gen6_block4_data(to_integer(unsigned(LUT_gen6_block4_addr)));
   LUT_gen6_block5_addr <= allbits(35 downto 30);
   LUT_gen6(5) <= LUT_gen6_block5_data(to_integer(unsigned(LUT_gen6_block5_addr)));
   LUT_gen6_block6_addr <= allbits(41 downto 36);
   LUT_gen6(6) <= LUT_gen6_block6_data(to_integer(unsigned(LUT_gen6_block6_addr)));
   LUT_gen6_block7_addr <= allbits(47 downto 42);
   LUT_gen6(7) <= LUT_gen6_block7_data(to_integer(unsigned(LUT_gen6_block7_addr)));
   LUT_gen6_block8_addr <= allbits(53 downto 48);
   LUT_gen6(8) <= LUT_gen6_block8_data(to_integer(unsigned(LUT_gen6_block8_addr)));
   LUT_gen6_block9_addr <= allbits(59 downto 54);
   LUT_gen6(9) <= LUT_gen6_block9_data(to_integer(unsigned(LUT_gen6_block9_addr)));
   LUT_gen6_block10_addr <= allbits(65 downto 60);
   LUT_gen6(10) <= LUT_gen6_block10_data(to_integer(unsigned(LUT_gen6_block10_addr)));
   LUT_gen6_block11_addr <= allbits(71 downto 66);
   LUT_gen6(11) <= LUT_gen6_block11_data(to_integer(unsigned(LUT_gen6_block11_addr)));
   LUT_gen6_block12_addr <= allbits(77 downto 72);
   LUT_gen6(12) <= LUT_gen6_block12_data(to_integer(unsigned(LUT_gen6_block12_addr)));
   LUT_gen6_block13_addr <= allbits(83 downto 78);
   LUT_gen6(13) <= LUT_gen6_block13_data(to_integer(unsigned(LUT_gen6_block13_addr)));
   LUT_gen6_block14_addr <= allbits(89 downto 84);
   LUT_gen6(14) <= LUT_gen6_block14_data(to_integer(unsigned(LUT_gen6_block14_addr)));
   LUT_gen6_block15_addr <= allbits(95 downto 90);
   LUT_gen6(15) <= LUT_gen6_block15_data(to_integer(unsigned(LUT_gen6_block15_addr)));
   LUT_gen7_block0_addr <= allbits(5 downto 0);
   LUT_gen7(0) <= LUT_gen7_block0_data(to_integer(unsigned(LUT_gen7_block0_addr)));
   LUT_gen7_block1_addr <= allbits(11 downto 6);
   LUT_gen7(1) <= LUT_gen7_block1_data(to_integer(unsigned(LUT_gen7_block1_addr)));
   LUT_gen7_block2_addr <= allbits(17 downto 12);
   LUT_gen7(2) <= LUT_gen7_block2_data(to_integer(unsigned(LUT_gen7_block2_addr)));
   LUT_gen7_block3_addr <= allbits(23 downto 18);
   LUT_gen7(3) <= LUT_gen7_block3_data(to_integer(unsigned(LUT_gen7_block3_addr)));
   LUT_gen7_block4_addr <= allbits(29 downto 24);
   LUT_gen7(4) <= LUT_gen7_block4_data(to_integer(unsigned(LUT_gen7_block4_addr)));
   LUT_gen7_block5_addr <= allbits(35 downto 30);
   LUT_gen7(5) <= LUT_gen7_block5_data(to_integer(unsigned(LUT_gen7_block5_addr)));
   LUT_gen7_block6_addr <= allbits(41 downto 36);
   LUT_gen7(6) <= LUT_gen7_block6_data(to_integer(unsigned(LUT_gen7_block6_addr)));
   LUT_gen7_block7_addr <= allbits(47 downto 42);
   LUT_gen7(7) <= LUT_gen7_block7_data(to_integer(unsigned(LUT_gen7_block7_addr)));
   LUT_gen7_block8_addr <= allbits(53 downto 48);
   LUT_gen7(8) <= LUT_gen7_block8_data(to_integer(unsigned(LUT_gen7_block8_addr)));
   LUT_gen7_block9_addr <= allbits(59 downto 54);
   LUT_gen7(9) <= LUT_gen7_block9_data(to_integer(unsigned(LUT_gen7_block9_addr)));
   LUT_gen7_block10_addr <= allbits(65 downto 60);
   LUT_gen7(10) <= LUT_gen7_block10_data(to_integer(unsigned(LUT_gen7_block10_addr)));
   LUT_gen7_block11_addr <= allbits(71 downto 66);
   LUT_gen7(11) <= LUT_gen7_block11_data(to_integer(unsigned(LUT_gen7_block11_addr)));
   LUT_gen7_block12_addr <= allbits(77 downto 72);
   LUT_gen7(12) <= LUT_gen7_block12_data(to_integer(unsigned(LUT_gen7_block12_addr)));
   LUT_gen7_block13_addr <= allbits(83 downto 78);
   LUT_gen7(13) <= LUT_gen7_block13_data(to_integer(unsigned(LUT_gen7_block13_addr)));
   LUT_gen7_block14_addr <= allbits(89 downto 84);
   LUT_gen7(14) <= LUT_gen7_block14_data(to_integer(unsigned(LUT_gen7_block14_addr)));
   LUT_gen7_block15_addr <= allbits(95 downto 90);
   LUT_gen7(15) <= LUT_gen7_block15_data(to_integer(unsigned(LUT_gen7_block15_addr)));
   LUT_gen8_block0_addr <= allbits(5 downto 0);
   LUT_gen8(0) <= LUT_gen8_block0_data(to_integer(unsigned(LUT_gen8_block0_addr)));
   LUT_gen8_block1_addr <= allbits(11 downto 6);
   LUT_gen8(1) <= LUT_gen8_block1_data(to_integer(unsigned(LUT_gen8_block1_addr)));
   LUT_gen8_block2_addr <= allbits(17 downto 12);
   LUT_gen8(2) <= LUT_gen8_block2_data(to_integer(unsigned(LUT_gen8_block2_addr)));
   LUT_gen8_block3_addr <= allbits(23 downto 18);
   LUT_gen8(3) <= LUT_gen8_block3_data(to_integer(unsigned(LUT_gen8_block3_addr)));
   LUT_gen8_block4_addr <= allbits(29 downto 24);
   LUT_gen8(4) <= LUT_gen8_block4_data(to_integer(unsigned(LUT_gen8_block4_addr)));
   LUT_gen8_block5_addr <= allbits(35 downto 30);
   LUT_gen8(5) <= LUT_gen8_block5_data(to_integer(unsigned(LUT_gen8_block5_addr)));
   LUT_gen8_block6_addr <= allbits(41 downto 36);
   LUT_gen8(6) <= LUT_gen8_block6_data(to_integer(unsigned(LUT_gen8_block6_addr)));
   LUT_gen8_block7_addr <= allbits(47 downto 42);
   LUT_gen8(7) <= LUT_gen8_block7_data(to_integer(unsigned(LUT_gen8_block7_addr)));
   LUT_gen8_block8_addr <= allbits(53 downto 48);
   LUT_gen8(8) <= LUT_gen8_block8_data(to_integer(unsigned(LUT_gen8_block8_addr)));
   LUT_gen8_block9_addr <= allbits(59 downto 54);
   LUT_gen8(9) <= LUT_gen8_block9_data(to_integer(unsigned(LUT_gen8_block9_addr)));
   LUT_gen8_block10_addr <= allbits(65 downto 60);
   LUT_gen8(10) <= LUT_gen8_block10_data(to_integer(unsigned(LUT_gen8_block10_addr)));
   LUT_gen8_block11_addr <= allbits(71 downto 66);
   LUT_gen8(11) <= LUT_gen8_block11_data(to_integer(unsigned(LUT_gen8_block11_addr)));
   LUT_gen8_block12_addr <= allbits(77 downto 72);
   LUT_gen8(12) <= LUT_gen8_block12_data(to_integer(unsigned(LUT_gen8_block12_addr)));
   LUT_gen8_block13_addr <= allbits(83 downto 78);
   LUT_gen8(13) <= LUT_gen8_block13_data(to_integer(unsigned(LUT_gen8_block13_addr)));
   LUT_gen8_block14_addr <= allbits(89 downto 84);
   LUT_gen8(14) <= LUT_gen8_block14_data(to_integer(unsigned(LUT_gen8_block14_addr)));
   LUT_gen8_block15_addr <= allbits(95 downto 90);
   LUT_gen8(15) <= LUT_gen8_block15_data(to_integer(unsigned(LUT_gen8_block15_addr)));
   LUT_gen9_block0_addr <= allbits(5 downto 0);
   LUT_gen9(0) <= LUT_gen9_block0_data(to_integer(unsigned(LUT_gen9_block0_addr)));
   LUT_gen9_block1_addr <= allbits(11 downto 6);
   LUT_gen9(1) <= LUT_gen9_block1_data(to_integer(unsigned(LUT_gen9_block1_addr)));
   LUT_gen9_block2_addr <= allbits(17 downto 12);
   LUT_gen9(2) <= LUT_gen9_block2_data(to_integer(unsigned(LUT_gen9_block2_addr)));
   LUT_gen9_block3_addr <= allbits(23 downto 18);
   LUT_gen9(3) <= LUT_gen9_block3_data(to_integer(unsigned(LUT_gen9_block3_addr)));
   LUT_gen9_block4_addr <= allbits(29 downto 24);
   LUT_gen9(4) <= LUT_gen9_block4_data(to_integer(unsigned(LUT_gen9_block4_addr)));
   LUT_gen9_block5_addr <= allbits(35 downto 30);
   LUT_gen9(5) <= LUT_gen9_block5_data(to_integer(unsigned(LUT_gen9_block5_addr)));
   LUT_gen9_block6_addr <= allbits(41 downto 36);
   LUT_gen9(6) <= LUT_gen9_block6_data(to_integer(unsigned(LUT_gen9_block6_addr)));
   LUT_gen9_block7_addr <= allbits(47 downto 42);
   LUT_gen9(7) <= LUT_gen9_block7_data(to_integer(unsigned(LUT_gen9_block7_addr)));
   LUT_gen9_block8_addr <= allbits(53 downto 48);
   LUT_gen9(8) <= LUT_gen9_block8_data(to_integer(unsigned(LUT_gen9_block8_addr)));
   LUT_gen9_block9_addr <= allbits(59 downto 54);
   LUT_gen9(9) <= LUT_gen9_block9_data(to_integer(unsigned(LUT_gen9_block9_addr)));
   LUT_gen9_block10_addr <= allbits(65 downto 60);
   LUT_gen9(10) <= LUT_gen9_block10_data(to_integer(unsigned(LUT_gen9_block10_addr)));
   LUT_gen9_block11_addr <= allbits(71 downto 66);
   LUT_gen9(11) <= LUT_gen9_block11_data(to_integer(unsigned(LUT_gen9_block11_addr)));
   LUT_gen9_block12_addr <= allbits(77 downto 72);
   LUT_gen9(12) <= LUT_gen9_block12_data(to_integer(unsigned(LUT_gen9_block12_addr)));
   LUT_gen9_block13_addr <= allbits(83 downto 78);
   LUT_gen9(13) <= LUT_gen9_block13_data(to_integer(unsigned(LUT_gen9_block13_addr)));
   LUT_gen9_block14_addr <= allbits(89 downto 84);
   LUT_gen9(14) <= LUT_gen9_block14_data(to_integer(unsigned(LUT_gen9_block14_addr)));
   LUT_gen9_block15_addr <= allbits(95 downto 90);
   LUT_gen9(15) <= LUT_gen9_block15_data(to_integer(unsigned(LUT_gen9_block15_addr)));
   LUT_gen10_block0_addr <= allbits(5 downto 0);
   LUT_gen10(0) <= LUT_gen10_block0_data(to_integer(unsigned(LUT_gen10_block0_addr)));
   LUT_gen10_block1_addr <= allbits(11 downto 6);
   LUT_gen10(1) <= LUT_gen10_block1_data(to_integer(unsigned(LUT_gen10_block1_addr)));
   LUT_gen10_block2_addr <= allbits(17 downto 12);
   LUT_gen10(2) <= LUT_gen10_block2_data(to_integer(unsigned(LUT_gen10_block2_addr)));
   LUT_gen10_block3_addr <= allbits(23 downto 18);
   LUT_gen10(3) <= LUT_gen10_block3_data(to_integer(unsigned(LUT_gen10_block3_addr)));
   LUT_gen10_block4_addr <= allbits(29 downto 24);
   LUT_gen10(4) <= LUT_gen10_block4_data(to_integer(unsigned(LUT_gen10_block4_addr)));
   LUT_gen10_block5_addr <= allbits(35 downto 30);
   LUT_gen10(5) <= LUT_gen10_block5_data(to_integer(unsigned(LUT_gen10_block5_addr)));
   LUT_gen10_block6_addr <= allbits(41 downto 36);
   LUT_gen10(6) <= LUT_gen10_block6_data(to_integer(unsigned(LUT_gen10_block6_addr)));
   LUT_gen10_block7_addr <= allbits(47 downto 42);
   LUT_gen10(7) <= LUT_gen10_block7_data(to_integer(unsigned(LUT_gen10_block7_addr)));
   LUT_gen10_block8_addr <= allbits(53 downto 48);
   LUT_gen10(8) <= LUT_gen10_block8_data(to_integer(unsigned(LUT_gen10_block8_addr)));
   LUT_gen10_block9_addr <= allbits(59 downto 54);
   LUT_gen10(9) <= LUT_gen10_block9_data(to_integer(unsigned(LUT_gen10_block9_addr)));
   LUT_gen10_block10_addr <= allbits(65 downto 60);
   LUT_gen10(10) <= LUT_gen10_block10_data(to_integer(unsigned(LUT_gen10_block10_addr)));
   LUT_gen10_block11_addr <= allbits(71 downto 66);
   LUT_gen10(11) <= LUT_gen10_block11_data(to_integer(unsigned(LUT_gen10_block11_addr)));
   LUT_gen10_block12_addr <= allbits(77 downto 72);
   LUT_gen10(12) <= LUT_gen10_block12_data(to_integer(unsigned(LUT_gen10_block12_addr)));
   LUT_gen10_block13_addr <= allbits(83 downto 78);
   LUT_gen10(13) <= LUT_gen10_block13_data(to_integer(unsigned(LUT_gen10_block13_addr)));
   LUT_gen10_block14_addr <= allbits(89 downto 84);
   LUT_gen10(14) <= LUT_gen10_block14_data(to_integer(unsigned(LUT_gen10_block14_addr)));
   LUT_gen10_block15_addr <= allbits(95 downto 90);
   LUT_gen10(15) <= LUT_gen10_block15_data(to_integer(unsigned(LUT_gen10_block15_addr)));
   LUT_gen11_block0_addr <= allbits(5 downto 0);
   LUT_gen11(0) <= LUT_gen11_block0_data(to_integer(unsigned(LUT_gen11_block0_addr)));
   LUT_gen11_block1_addr <= allbits(11 downto 6);
   LUT_gen11(1) <= LUT_gen11_block1_data(to_integer(unsigned(LUT_gen11_block1_addr)));
   LUT_gen11_block2_addr <= allbits(17 downto 12);
   LUT_gen11(2) <= LUT_gen11_block2_data(to_integer(unsigned(LUT_gen11_block2_addr)));
   LUT_gen11_block3_addr <= allbits(23 downto 18);
   LUT_gen11(3) <= LUT_gen11_block3_data(to_integer(unsigned(LUT_gen11_block3_addr)));
   LUT_gen11_block4_addr <= allbits(29 downto 24);
   LUT_gen11(4) <= LUT_gen11_block4_data(to_integer(unsigned(LUT_gen11_block4_addr)));
   LUT_gen11_block5_addr <= allbits(35 downto 30);
   LUT_gen11(5) <= LUT_gen11_block5_data(to_integer(unsigned(LUT_gen11_block5_addr)));
   LUT_gen11_block6_addr <= allbits(41 downto 36);
   LUT_gen11(6) <= LUT_gen11_block6_data(to_integer(unsigned(LUT_gen11_block6_addr)));
   LUT_gen11_block7_addr <= allbits(47 downto 42);
   LUT_gen11(7) <= LUT_gen11_block7_data(to_integer(unsigned(LUT_gen11_block7_addr)));
   LUT_gen11(8) <= '0';
   LUT_gen11_block9_addr <= allbits(59 downto 54);
   LUT_gen11(9) <= LUT_gen11_block9_data(to_integer(unsigned(LUT_gen11_block9_addr)));
   LUT_gen11_block10_addr <= allbits(65 downto 60);
   LUT_gen11(10) <= LUT_gen11_block10_data(to_integer(unsigned(LUT_gen11_block10_addr)));
   LUT_gen11_block11_addr <= allbits(71 downto 66);
   LUT_gen11(11) <= LUT_gen11_block11_data(to_integer(unsigned(LUT_gen11_block11_addr)));
   LUT_gen11_block12_addr <= allbits(77 downto 72);
   LUT_gen11(12) <= LUT_gen11_block12_data(to_integer(unsigned(LUT_gen11_block12_addr)));
   LUT_gen11_block13_addr <= allbits(83 downto 78);
   LUT_gen11(13) <= LUT_gen11_block13_data(to_integer(unsigned(LUT_gen11_block13_addr)));
   LUT_gen11_block14_addr <= allbits(89 downto 84);
   LUT_gen11(14) <= LUT_gen11_block14_data(to_integer(unsigned(LUT_gen11_block14_addr)));
   LUT_gen11_block15_addr <= allbits(95 downto 90);
   LUT_gen11(15) <= LUT_gen11_block15_data(to_integer(unsigned(LUT_gen11_block15_addr)));
   LUT_gen12_block0_addr <= allbits(5 downto 0);
   LUT_gen12(0) <= LUT_gen12_block0_data(to_integer(unsigned(LUT_gen12_block0_addr)));
   LUT_gen12_block1_addr <= allbits(11 downto 6);
   LUT_gen12(1) <= LUT_gen12_block1_data(to_integer(unsigned(LUT_gen12_block1_addr)));
   LUT_gen12_block2_addr <= allbits(17 downto 12);
   LUT_gen12(2) <= LUT_gen12_block2_data(to_integer(unsigned(LUT_gen12_block2_addr)));
   LUT_gen12_block3_addr <= allbits(23 downto 18);
   LUT_gen12(3) <= LUT_gen12_block3_data(to_integer(unsigned(LUT_gen12_block3_addr)));
   LUT_gen12_block4_addr <= allbits(29 downto 24);
   LUT_gen12(4) <= LUT_gen12_block4_data(to_integer(unsigned(LUT_gen12_block4_addr)));
   LUT_gen12_block5_addr <= allbits(35 downto 30);
   LUT_gen12(5) <= LUT_gen12_block5_data(to_integer(unsigned(LUT_gen12_block5_addr)));
   LUT_gen12_block6_addr <= allbits(41 downto 36);
   LUT_gen12(6) <= LUT_gen12_block6_data(to_integer(unsigned(LUT_gen12_block6_addr)));
   LUT_gen12_block7_addr <= allbits(47 downto 42);
   LUT_gen12(7) <= LUT_gen12_block7_data(to_integer(unsigned(LUT_gen12_block7_addr)));
   LUT_gen12_block8_addr <= allbits(53 downto 48);
   LUT_gen12(8) <= LUT_gen12_block8_data(to_integer(unsigned(LUT_gen12_block8_addr)));
   LUT_gen12_block9_addr <= allbits(59 downto 54);
   LUT_gen12(9) <= LUT_gen12_block9_data(to_integer(unsigned(LUT_gen12_block9_addr)));
   LUT_gen12_block10_addr <= allbits(65 downto 60);
   LUT_gen12(10) <= LUT_gen12_block10_data(to_integer(unsigned(LUT_gen12_block10_addr)));
   LUT_gen12_block11_addr <= allbits(71 downto 66);
   LUT_gen12(11) <= LUT_gen12_block11_data(to_integer(unsigned(LUT_gen12_block11_addr)));
   LUT_gen12_block12_addr <= allbits(77 downto 72);
   LUT_gen12(12) <= LUT_gen12_block12_data(to_integer(unsigned(LUT_gen12_block12_addr)));
   LUT_gen12_block13_addr <= allbits(83 downto 78);
   LUT_gen12(13) <= LUT_gen12_block13_data(to_integer(unsigned(LUT_gen12_block13_addr)));
   LUT_gen12_block14_addr <= allbits(89 downto 84);
   LUT_gen12(14) <= LUT_gen12_block14_data(to_integer(unsigned(LUT_gen12_block14_addr)));
   LUT_gen12_block15_addr <= allbits(95 downto 90);
   LUT_gen12(15) <= LUT_gen12_block15_data(to_integer(unsigned(LUT_gen12_block15_addr)));
   LUT_gen13_block0_addr <= allbits(5 downto 0);
   LUT_gen13(0) <= LUT_gen13_block0_data(to_integer(unsigned(LUT_gen13_block0_addr)));
   LUT_gen13_block1_addr <= allbits(11 downto 6);
   LUT_gen13(1) <= LUT_gen13_block1_data(to_integer(unsigned(LUT_gen13_block1_addr)));
   LUT_gen13_block2_addr <= allbits(17 downto 12);
   LUT_gen13(2) <= LUT_gen13_block2_data(to_integer(unsigned(LUT_gen13_block2_addr)));
   LUT_gen13(3) <= '0';
   LUT_gen13_block4_addr <= allbits(29 downto 24);
   LUT_gen13(4) <= LUT_gen13_block4_data(to_integer(unsigned(LUT_gen13_block4_addr)));
   LUT_gen13_block5_addr <= allbits(35 downto 30);
   LUT_gen13(5) <= LUT_gen13_block5_data(to_integer(unsigned(LUT_gen13_block5_addr)));
   LUT_gen13_block6_addr <= allbits(41 downto 36);
   LUT_gen13(6) <= LUT_gen13_block6_data(to_integer(unsigned(LUT_gen13_block6_addr)));
   LUT_gen13_block7_addr <= allbits(47 downto 42);
   LUT_gen13(7) <= LUT_gen13_block7_data(to_integer(unsigned(LUT_gen13_block7_addr)));
   LUT_gen13_block8_addr <= allbits(53 downto 48);
   LUT_gen13(8) <= LUT_gen13_block8_data(to_integer(unsigned(LUT_gen13_block8_addr)));
   LUT_gen13_block9_addr <= allbits(59 downto 54);
   LUT_gen13(9) <= LUT_gen13_block9_data(to_integer(unsigned(LUT_gen13_block9_addr)));
   LUT_gen13_block10_addr <= allbits(65 downto 60);
   LUT_gen13(10) <= LUT_gen13_block10_data(to_integer(unsigned(LUT_gen13_block10_addr)));
   LUT_gen13_block11_addr <= allbits(71 downto 66);
   LUT_gen13(11) <= LUT_gen13_block11_data(to_integer(unsigned(LUT_gen13_block11_addr)));
   LUT_gen13_block12_addr <= allbits(77 downto 72);
   LUT_gen13(12) <= LUT_gen13_block12_data(to_integer(unsigned(LUT_gen13_block12_addr)));
   LUT_gen13_block13_addr <= allbits(83 downto 78);
   LUT_gen13(13) <= LUT_gen13_block13_data(to_integer(unsigned(LUT_gen13_block13_addr)));
   LUT_gen13_block14_addr <= allbits(89 downto 84);
   LUT_gen13(14) <= LUT_gen13_block14_data(to_integer(unsigned(LUT_gen13_block14_addr)));
   LUT_gen13_block15_addr <= allbits(95 downto 90);
   LUT_gen13(15) <= LUT_gen13_block15_data(to_integer(unsigned(LUT_gen13_block15_addr)));
   LUT_gen14_block0_addr <= allbits(5 downto 0);
   LUT_gen14(0) <= LUT_gen14_block0_data(to_integer(unsigned(LUT_gen14_block0_addr)));
   LUT_gen14_block1_addr <= allbits(11 downto 6);
   LUT_gen14(1) <= LUT_gen14_block1_data(to_integer(unsigned(LUT_gen14_block1_addr)));
   LUT_gen14_block2_addr <= allbits(17 downto 12);
   LUT_gen14(2) <= LUT_gen14_block2_data(to_integer(unsigned(LUT_gen14_block2_addr)));
   LUT_gen14_block3_addr <= allbits(23 downto 18);
   LUT_gen14(3) <= LUT_gen14_block3_data(to_integer(unsigned(LUT_gen14_block3_addr)));
   LUT_gen14_block4_addr <= allbits(29 downto 24);
   LUT_gen14(4) <= LUT_gen14_block4_data(to_integer(unsigned(LUT_gen14_block4_addr)));
   LUT_gen14_block5_addr <= allbits(35 downto 30);
   LUT_gen14(5) <= LUT_gen14_block5_data(to_integer(unsigned(LUT_gen14_block5_addr)));
   LUT_gen14_block6_addr <= allbits(41 downto 36);
   LUT_gen14(6) <= LUT_gen14_block6_data(to_integer(unsigned(LUT_gen14_block6_addr)));
   LUT_gen14_block7_addr <= allbits(47 downto 42);
   LUT_gen14(7) <= LUT_gen14_block7_data(to_integer(unsigned(LUT_gen14_block7_addr)));
   LUT_gen14_block8_addr <= allbits(53 downto 48);
   LUT_gen14(8) <= LUT_gen14_block8_data(to_integer(unsigned(LUT_gen14_block8_addr)));
   LUT_gen14_block9_addr <= allbits(59 downto 54);
   LUT_gen14(9) <= LUT_gen14_block9_data(to_integer(unsigned(LUT_gen14_block9_addr)));
   LUT_gen14_block10_addr <= allbits(65 downto 60);
   LUT_gen14(10) <= LUT_gen14_block10_data(to_integer(unsigned(LUT_gen14_block10_addr)));
   LUT_gen14_block11_addr <= allbits(71 downto 66);
   LUT_gen14(11) <= LUT_gen14_block11_data(to_integer(unsigned(LUT_gen14_block11_addr)));
   LUT_gen14_block12_addr <= allbits(77 downto 72);
   LUT_gen14(12) <= LUT_gen14_block12_data(to_integer(unsigned(LUT_gen14_block12_addr)));
   LUT_gen14_block13_addr <= allbits(83 downto 78);
   LUT_gen14(13) <= LUT_gen14_block13_data(to_integer(unsigned(LUT_gen14_block13_addr)));
   LUT_gen14_block14_addr <= allbits(89 downto 84);
   LUT_gen14(14) <= LUT_gen14_block14_data(to_integer(unsigned(LUT_gen14_block14_addr)));
   LUT_gen14_block15_addr <= allbits(95 downto 90);
   LUT_gen14(15) <= LUT_gen14_block15_data(to_integer(unsigned(LUT_gen14_block15_addr)));
   LUT_gen15(0) <= '0';
   LUT_gen15_block1_addr <= allbits(11 downto 6);
   LUT_gen15(1) <= LUT_gen15_block1_data(to_integer(unsigned(LUT_gen15_block1_addr)));
   LUT_gen15_block2_addr <= allbits(17 downto 12);
   LUT_gen15(2) <= LUT_gen15_block2_data(to_integer(unsigned(LUT_gen15_block2_addr)));
   LUT_gen15_block3_addr <= allbits(23 downto 18);
   LUT_gen15(3) <= LUT_gen15_block3_data(to_integer(unsigned(LUT_gen15_block3_addr)));
   LUT_gen15_block4_addr <= allbits(29 downto 24);
   LUT_gen15(4) <= LUT_gen15_block4_data(to_integer(unsigned(LUT_gen15_block4_addr)));
   LUT_gen15_block5_addr <= allbits(35 downto 30);
   LUT_gen15(5) <= LUT_gen15_block5_data(to_integer(unsigned(LUT_gen15_block5_addr)));
   LUT_gen15_block6_addr <= allbits(41 downto 36);
   LUT_gen15(6) <= LUT_gen15_block6_data(to_integer(unsigned(LUT_gen15_block6_addr)));
   LUT_gen15_block7_addr <= allbits(47 downto 42);
   LUT_gen15(7) <= LUT_gen15_block7_data(to_integer(unsigned(LUT_gen15_block7_addr)));
   LUT_gen15_block8_addr <= allbits(53 downto 48);
   LUT_gen15(8) <= LUT_gen15_block8_data(to_integer(unsigned(LUT_gen15_block8_addr)));
   LUT_gen15_block9_addr <= allbits(59 downto 54);
   LUT_gen15(9) <= LUT_gen15_block9_data(to_integer(unsigned(LUT_gen15_block9_addr)));
   LUT_gen15_block10_addr <= allbits(65 downto 60);
   LUT_gen15(10) <= LUT_gen15_block10_data(to_integer(unsigned(LUT_gen15_block10_addr)));
   LUT_gen15_block11_addr <= allbits(71 downto 66);
   LUT_gen15(11) <= LUT_gen15_block11_data(to_integer(unsigned(LUT_gen15_block11_addr)));
   LUT_gen15_block12_addr <= allbits(77 downto 72);
   LUT_gen15(12) <= LUT_gen15_block12_data(to_integer(unsigned(LUT_gen15_block12_addr)));
   LUT_gen15_block13_addr <= allbits(83 downto 78);
   LUT_gen15(13) <= LUT_gen15_block13_data(to_integer(unsigned(LUT_gen15_block13_addr)));
   LUT_gen15_block14_addr <= allbits(89 downto 84);
   LUT_gen15(14) <= LUT_gen15_block14_data(to_integer(unsigned(LUT_gen15_block14_addr)));
   LUT_gen15_block15_addr <= allbits(95 downto 90);
   LUT_gen15(15) <= LUT_gen15_block15_data(to_integer(unsigned(LUT_gen15_block15_addr)));
   LUT_gen16_block0_addr <= allbits(5 downto 0);
   LUT_gen16(0) <= LUT_gen16_block0_data(to_integer(unsigned(LUT_gen16_block0_addr)));
   LUT_gen16_block1_addr <= allbits(11 downto 6);
   LUT_gen16(1) <= LUT_gen16_block1_data(to_integer(unsigned(LUT_gen16_block1_addr)));
   LUT_gen16_block2_addr <= allbits(17 downto 12);
   LUT_gen16(2) <= LUT_gen16_block2_data(to_integer(unsigned(LUT_gen16_block2_addr)));
   LUT_gen16_block3_addr <= allbits(23 downto 18);
   LUT_gen16(3) <= LUT_gen16_block3_data(to_integer(unsigned(LUT_gen16_block3_addr)));
   LUT_gen16_block4_addr <= allbits(29 downto 24);
   LUT_gen16(4) <= LUT_gen16_block4_data(to_integer(unsigned(LUT_gen16_block4_addr)));
   LUT_gen16_block5_addr <= allbits(35 downto 30);
   LUT_gen16(5) <= LUT_gen16_block5_data(to_integer(unsigned(LUT_gen16_block5_addr)));
   LUT_gen16_block6_addr <= allbits(41 downto 36);
   LUT_gen16(6) <= LUT_gen16_block6_data(to_integer(unsigned(LUT_gen16_block6_addr)));
   LUT_gen16_block7_addr <= allbits(47 downto 42);
   LUT_gen16(7) <= LUT_gen16_block7_data(to_integer(unsigned(LUT_gen16_block7_addr)));
   LUT_gen16_block8_addr <= allbits(53 downto 48);
   LUT_gen16(8) <= LUT_gen16_block8_data(to_integer(unsigned(LUT_gen16_block8_addr)));
   LUT_gen16(9) <= '0';
   LUT_gen16_block10_addr <= allbits(65 downto 60);
   LUT_gen16(10) <= LUT_gen16_block10_data(to_integer(unsigned(LUT_gen16_block10_addr)));
   LUT_gen16_block11_addr <= allbits(71 downto 66);
   LUT_gen16(11) <= LUT_gen16_block11_data(to_integer(unsigned(LUT_gen16_block11_addr)));
   LUT_gen16_block12_addr <= allbits(77 downto 72);
   LUT_gen16(12) <= LUT_gen16_block12_data(to_integer(unsigned(LUT_gen16_block12_addr)));
   LUT_gen16_block13_addr <= allbits(83 downto 78);
   LUT_gen16(13) <= LUT_gen16_block13_data(to_integer(unsigned(LUT_gen16_block13_addr)));
   LUT_gen16_block14_addr <= allbits(89 downto 84);
   LUT_gen16(14) <= LUT_gen16_block14_data(to_integer(unsigned(LUT_gen16_block14_addr)));
   LUT_gen16_block15_addr <= allbits(95 downto 90);
   LUT_gen16(15) <= LUT_gen16_block15_data(to_integer(unsigned(LUT_gen16_block15_addr)));
   LUT_gen17_block0_addr <= allbits(5 downto 0);
   LUT_gen17(0) <= LUT_gen17_block0_data(to_integer(unsigned(LUT_gen17_block0_addr)));
   LUT_gen17_block1_addr <= allbits(11 downto 6);
   LUT_gen17(1) <= LUT_gen17_block1_data(to_integer(unsigned(LUT_gen17_block1_addr)));
   LUT_gen17_block2_addr <= allbits(17 downto 12);
   LUT_gen17(2) <= LUT_gen17_block2_data(to_integer(unsigned(LUT_gen17_block2_addr)));
   LUT_gen17_block3_addr <= allbits(23 downto 18);
   LUT_gen17(3) <= LUT_gen17_block3_data(to_integer(unsigned(LUT_gen17_block3_addr)));
   LUT_gen17(4) <= '0';
   LUT_gen17_block5_addr <= allbits(35 downto 30);
   LUT_gen17(5) <= LUT_gen17_block5_data(to_integer(unsigned(LUT_gen17_block5_addr)));
   LUT_gen17_block6_addr <= allbits(41 downto 36);
   LUT_gen17(6) <= LUT_gen17_block6_data(to_integer(unsigned(LUT_gen17_block6_addr)));
   LUT_gen17_block7_addr <= allbits(47 downto 42);
   LUT_gen17(7) <= LUT_gen17_block7_data(to_integer(unsigned(LUT_gen17_block7_addr)));
   LUT_gen17_block8_addr <= allbits(53 downto 48);
   LUT_gen17(8) <= LUT_gen17_block8_data(to_integer(unsigned(LUT_gen17_block8_addr)));
   LUT_gen17(9) <= '0';
   LUT_gen17_block10_addr <= allbits(65 downto 60);
   LUT_gen17(10) <= LUT_gen17_block10_data(to_integer(unsigned(LUT_gen17_block10_addr)));
   LUT_gen17_block11_addr <= allbits(71 downto 66);
   LUT_gen17(11) <= LUT_gen17_block11_data(to_integer(unsigned(LUT_gen17_block11_addr)));
   LUT_gen17_block12_addr <= allbits(77 downto 72);
   LUT_gen17(12) <= LUT_gen17_block12_data(to_integer(unsigned(LUT_gen17_block12_addr)));
   LUT_gen17_block13_addr <= allbits(83 downto 78);
   LUT_gen17(13) <= LUT_gen17_block13_data(to_integer(unsigned(LUT_gen17_block13_addr)));
   LUT_gen17_block14_addr <= allbits(89 downto 84);
   LUT_gen17(14) <= LUT_gen17_block14_data(to_integer(unsigned(LUT_gen17_block14_addr)));
   LUT_gen17_block15_addr <= allbits(95 downto 90);
   LUT_gen17(15) <= LUT_gen17_block15_data(to_integer(unsigned(LUT_gen17_block15_addr)));
   LUT_gen18_block0_addr <= allbits(5 downto 0);
   LUT_gen18(0) <= LUT_gen18_block0_data(to_integer(unsigned(LUT_gen18_block0_addr)));
   LUT_gen18_block1_addr <= allbits(11 downto 6);
   LUT_gen18(1) <= LUT_gen18_block1_data(to_integer(unsigned(LUT_gen18_block1_addr)));
   LUT_gen18_block2_addr <= allbits(17 downto 12);
   LUT_gen18(2) <= LUT_gen18_block2_data(to_integer(unsigned(LUT_gen18_block2_addr)));
   LUT_gen18_block3_addr <= allbits(23 downto 18);
   LUT_gen18(3) <= LUT_gen18_block3_data(to_integer(unsigned(LUT_gen18_block3_addr)));
   LUT_gen18(4) <= '0';
   LUT_gen18_block5_addr <= allbits(35 downto 30);
   LUT_gen18(5) <= LUT_gen18_block5_data(to_integer(unsigned(LUT_gen18_block5_addr)));
   LUT_gen18_block6_addr <= allbits(41 downto 36);
   LUT_gen18(6) <= LUT_gen18_block6_data(to_integer(unsigned(LUT_gen18_block6_addr)));
   LUT_gen18_block7_addr <= allbits(47 downto 42);
   LUT_gen18(7) <= LUT_gen18_block7_data(to_integer(unsigned(LUT_gen18_block7_addr)));
   LUT_gen18_block8_addr <= allbits(53 downto 48);
   LUT_gen18(8) <= LUT_gen18_block8_data(to_integer(unsigned(LUT_gen18_block8_addr)));
   LUT_gen18(9) <= '0';
   LUT_gen18_block10_addr <= allbits(65 downto 60);
   LUT_gen18(10) <= LUT_gen18_block10_data(to_integer(unsigned(LUT_gen18_block10_addr)));
   LUT_gen18_block11_addr <= allbits(71 downto 66);
   LUT_gen18(11) <= LUT_gen18_block11_data(to_integer(unsigned(LUT_gen18_block11_addr)));
   LUT_gen18_block12_addr <= allbits(77 downto 72);
   LUT_gen18(12) <= LUT_gen18_block12_data(to_integer(unsigned(LUT_gen18_block12_addr)));
   LUT_gen18_block13_addr <= allbits(83 downto 78);
   LUT_gen18(13) <= LUT_gen18_block13_data(to_integer(unsigned(LUT_gen18_block13_addr)));
   LUT_gen18_block14_addr <= allbits(89 downto 84);
   LUT_gen18(14) <= LUT_gen18_block14_data(to_integer(unsigned(LUT_gen18_block14_addr)));
   LUT_gen18_block15_addr <= allbits(95 downto 90);
   LUT_gen18(15) <= LUT_gen18_block15_data(to_integer(unsigned(LUT_gen18_block15_addr)));
   LUT_gen19_block0_addr <= allbits(5 downto 0);
   LUT_gen19(0) <= LUT_gen19_block0_data(to_integer(unsigned(LUT_gen19_block0_addr)));
   LUT_gen19_block1_addr <= allbits(11 downto 6);
   LUT_gen19(1) <= LUT_gen19_block1_data(to_integer(unsigned(LUT_gen19_block1_addr)));
   LUT_gen19_block2_addr <= allbits(17 downto 12);
   LUT_gen19(2) <= LUT_gen19_block2_data(to_integer(unsigned(LUT_gen19_block2_addr)));
   LUT_gen19_block3_addr <= allbits(23 downto 18);
   LUT_gen19(3) <= LUT_gen19_block3_data(to_integer(unsigned(LUT_gen19_block3_addr)));
   LUT_gen19(4) <= '0';
   LUT_gen19_block5_addr <= allbits(35 downto 30);
   LUT_gen19(5) <= LUT_gen19_block5_data(to_integer(unsigned(LUT_gen19_block5_addr)));
   LUT_gen19_block6_addr <= allbits(41 downto 36);
   LUT_gen19(6) <= LUT_gen19_block6_data(to_integer(unsigned(LUT_gen19_block6_addr)));
   LUT_gen19_block7_addr <= allbits(47 downto 42);
   LUT_gen19(7) <= LUT_gen19_block7_data(to_integer(unsigned(LUT_gen19_block7_addr)));
   LUT_gen19_block8_addr <= allbits(53 downto 48);
   LUT_gen19(8) <= LUT_gen19_block8_data(to_integer(unsigned(LUT_gen19_block8_addr)));
   LUT_gen19_block9_addr <= allbits(59 downto 54);
   LUT_gen19(9) <= LUT_gen19_block9_data(to_integer(unsigned(LUT_gen19_block9_addr)));
   LUT_gen19_block10_addr <= allbits(65 downto 60);
   LUT_gen19(10) <= LUT_gen19_block10_data(to_integer(unsigned(LUT_gen19_block10_addr)));
   LUT_gen19_block11_addr <= allbits(71 downto 66);
   LUT_gen19(11) <= LUT_gen19_block11_data(to_integer(unsigned(LUT_gen19_block11_addr)));
   LUT_gen19_block12_addr <= allbits(77 downto 72);
   LUT_gen19(12) <= LUT_gen19_block12_data(to_integer(unsigned(LUT_gen19_block12_addr)));
   LUT_gen19_block13_addr <= allbits(83 downto 78);
   LUT_gen19(13) <= LUT_gen19_block13_data(to_integer(unsigned(LUT_gen19_block13_addr)));
   LUT_gen19_block14_addr <= allbits(89 downto 84);
   LUT_gen19(14) <= LUT_gen19_block14_data(to_integer(unsigned(LUT_gen19_block14_addr)));
   LUT_gen19_block15_addr <= allbits(95 downto 90);
   LUT_gen19(15) <= LUT_gen19_block15_data(to_integer(unsigned(LUT_gen19_block15_addr)));
   LUT_gen20_block0_addr <= allbits(5 downto 0);
   LUT_gen20(0) <= LUT_gen20_block0_data(to_integer(unsigned(LUT_gen20_block0_addr)));
   LUT_gen20_block1_addr <= allbits(11 downto 6);
   LUT_gen20(1) <= LUT_gen20_block1_data(to_integer(unsigned(LUT_gen20_block1_addr)));
   LUT_gen20_block2_addr <= allbits(17 downto 12);
   LUT_gen20(2) <= LUT_gen20_block2_data(to_integer(unsigned(LUT_gen20_block2_addr)));
   LUT_gen20_block3_addr <= allbits(23 downto 18);
   LUT_gen20(3) <= LUT_gen20_block3_data(to_integer(unsigned(LUT_gen20_block3_addr)));
   LUT_gen20_block4_addr <= allbits(29 downto 24);
   LUT_gen20(4) <= LUT_gen20_block4_data(to_integer(unsigned(LUT_gen20_block4_addr)));
   LUT_gen20_block5_addr <= allbits(35 downto 30);
   LUT_gen20(5) <= LUT_gen20_block5_data(to_integer(unsigned(LUT_gen20_block5_addr)));
   LUT_gen20_block6_addr <= allbits(41 downto 36);
   LUT_gen20(6) <= LUT_gen20_block6_data(to_integer(unsigned(LUT_gen20_block6_addr)));
   LUT_gen20_block7_addr <= allbits(47 downto 42);
   LUT_gen20(7) <= LUT_gen20_block7_data(to_integer(unsigned(LUT_gen20_block7_addr)));
   LUT_gen20_block8_addr <= allbits(53 downto 48);
   LUT_gen20(8) <= LUT_gen20_block8_data(to_integer(unsigned(LUT_gen20_block8_addr)));
   LUT_gen20_block9_addr <= allbits(59 downto 54);
   LUT_gen20(9) <= LUT_gen20_block9_data(to_integer(unsigned(LUT_gen20_block9_addr)));
   LUT_gen20_block10_addr <= allbits(65 downto 60);
   LUT_gen20(10) <= LUT_gen20_block10_data(to_integer(unsigned(LUT_gen20_block10_addr)));
   LUT_gen20_block11_addr <= allbits(71 downto 66);
   LUT_gen20(11) <= LUT_gen20_block11_data(to_integer(unsigned(LUT_gen20_block11_addr)));
   LUT_gen20_block12_addr <= allbits(77 downto 72);
   LUT_gen20(12) <= LUT_gen20_block12_data(to_integer(unsigned(LUT_gen20_block12_addr)));
   LUT_gen20_block13_addr <= allbits(83 downto 78);
   LUT_gen20(13) <= LUT_gen20_block13_data(to_integer(unsigned(LUT_gen20_block13_addr)));
   LUT_gen20_block14_addr <= allbits(89 downto 84);
   LUT_gen20(14) <= LUT_gen20_block14_data(to_integer(unsigned(LUT_gen20_block14_addr)));
   LUT_gen20_block15_addr <= allbits(95 downto 90);
   LUT_gen20(15) <= LUT_gen20_block15_data(to_integer(unsigned(LUT_gen20_block15_addr)));
   LUT_gen21_block0_addr <= allbits(5 downto 0);
   LUT_gen21(0) <= LUT_gen21_block0_data(to_integer(unsigned(LUT_gen21_block0_addr)));
   LUT_gen21_block1_addr <= allbits(11 downto 6);
   LUT_gen21(1) <= LUT_gen21_block1_data(to_integer(unsigned(LUT_gen21_block1_addr)));
   LUT_gen21_block2_addr <= allbits(17 downto 12);
   LUT_gen21(2) <= LUT_gen21_block2_data(to_integer(unsigned(LUT_gen21_block2_addr)));
   LUT_gen21_block3_addr <= allbits(23 downto 18);
   LUT_gen21(3) <= LUT_gen21_block3_data(to_integer(unsigned(LUT_gen21_block3_addr)));
   LUT_gen21_block4_addr <= allbits(29 downto 24);
   LUT_gen21(4) <= LUT_gen21_block4_data(to_integer(unsigned(LUT_gen21_block4_addr)));
   LUT_gen21_block5_addr <= allbits(35 downto 30);
   LUT_gen21(5) <= LUT_gen21_block5_data(to_integer(unsigned(LUT_gen21_block5_addr)));
   LUT_gen21_block6_addr <= allbits(41 downto 36);
   LUT_gen21(6) <= LUT_gen21_block6_data(to_integer(unsigned(LUT_gen21_block6_addr)));
   LUT_gen21_block7_addr <= allbits(47 downto 42);
   LUT_gen21(7) <= LUT_gen21_block7_data(to_integer(unsigned(LUT_gen21_block7_addr)));
   LUT_gen21_block8_addr <= allbits(53 downto 48);
   LUT_gen21(8) <= LUT_gen21_block8_data(to_integer(unsigned(LUT_gen21_block8_addr)));
   LUT_gen21_block9_addr <= allbits(59 downto 54);
   LUT_gen21(9) <= LUT_gen21_block9_data(to_integer(unsigned(LUT_gen21_block9_addr)));
   LUT_gen21_block10_addr <= allbits(65 downto 60);
   LUT_gen21(10) <= LUT_gen21_block10_data(to_integer(unsigned(LUT_gen21_block10_addr)));
   LUT_gen21_block11_addr <= allbits(71 downto 66);
   LUT_gen21(11) <= LUT_gen21_block11_data(to_integer(unsigned(LUT_gen21_block11_addr)));
   LUT_gen21_block12_addr <= allbits(77 downto 72);
   LUT_gen21(12) <= LUT_gen21_block12_data(to_integer(unsigned(LUT_gen21_block12_addr)));
   LUT_gen21_block13_addr <= allbits(83 downto 78);
   LUT_gen21(13) <= LUT_gen21_block13_data(to_integer(unsigned(LUT_gen21_block13_addr)));
   LUT_gen21_block14_addr <= allbits(89 downto 84);
   LUT_gen21(14) <= LUT_gen21_block14_data(to_integer(unsigned(LUT_gen21_block14_addr)));
   LUT_gen21_block15_addr <= allbits(95 downto 90);
   LUT_gen21(15) <= LUT_gen21_block15_data(to_integer(unsigned(LUT_gen21_block15_addr)));
   LUT_gen22_block0_addr <= allbits(5 downto 0);
   LUT_gen22(0) <= LUT_gen22_block0_data(to_integer(unsigned(LUT_gen22_block0_addr)));
   LUT_gen22_block1_addr <= allbits(11 downto 6);
   LUT_gen22(1) <= LUT_gen22_block1_data(to_integer(unsigned(LUT_gen22_block1_addr)));
   LUT_gen22_block2_addr <= allbits(17 downto 12);
   LUT_gen22(2) <= LUT_gen22_block2_data(to_integer(unsigned(LUT_gen22_block2_addr)));
   LUT_gen22_block3_addr <= allbits(23 downto 18);
   LUT_gen22(3) <= LUT_gen22_block3_data(to_integer(unsigned(LUT_gen22_block3_addr)));
   LUT_gen22_block4_addr <= allbits(29 downto 24);
   LUT_gen22(4) <= LUT_gen22_block4_data(to_integer(unsigned(LUT_gen22_block4_addr)));
   LUT_gen22_block5_addr <= allbits(35 downto 30);
   LUT_gen22(5) <= LUT_gen22_block5_data(to_integer(unsigned(LUT_gen22_block5_addr)));
   LUT_gen22_block6_addr <= allbits(41 downto 36);
   LUT_gen22(6) <= LUT_gen22_block6_data(to_integer(unsigned(LUT_gen22_block6_addr)));
   LUT_gen22_block7_addr <= allbits(47 downto 42);
   LUT_gen22(7) <= LUT_gen22_block7_data(to_integer(unsigned(LUT_gen22_block7_addr)));
   LUT_gen22_block8_addr <= allbits(53 downto 48);
   LUT_gen22(8) <= LUT_gen22_block8_data(to_integer(unsigned(LUT_gen22_block8_addr)));
   LUT_gen22_block9_addr <= allbits(59 downto 54);
   LUT_gen22(9) <= LUT_gen22_block9_data(to_integer(unsigned(LUT_gen22_block9_addr)));
   LUT_gen22_block10_addr <= allbits(65 downto 60);
   LUT_gen22(10) <= LUT_gen22_block10_data(to_integer(unsigned(LUT_gen22_block10_addr)));
   LUT_gen22_block11_addr <= allbits(71 downto 66);
   LUT_gen22(11) <= LUT_gen22_block11_data(to_integer(unsigned(LUT_gen22_block11_addr)));
   LUT_gen22_block12_addr <= allbits(77 downto 72);
   LUT_gen22(12) <= LUT_gen22_block12_data(to_integer(unsigned(LUT_gen22_block12_addr)));
   LUT_gen22_block13_addr <= allbits(83 downto 78);
   LUT_gen22(13) <= LUT_gen22_block13_data(to_integer(unsigned(LUT_gen22_block13_addr)));
   LUT_gen22_block14_addr <= allbits(89 downto 84);
   LUT_gen22(14) <= LUT_gen22_block14_data(to_integer(unsigned(LUT_gen22_block14_addr)));
   LUT_gen22_block15_addr <= allbits(95 downto 90);
   LUT_gen22(15) <= LUT_gen22_block15_data(to_integer(unsigned(LUT_gen22_block15_addr)));
   LUT_gen23_block0_addr <= allbits(5 downto 0);
   LUT_gen23(0) <= LUT_gen23_block0_data(to_integer(unsigned(LUT_gen23_block0_addr)));
   LUT_gen23_block1_addr <= allbits(11 downto 6);
   LUT_gen23(1) <= LUT_gen23_block1_data(to_integer(unsigned(LUT_gen23_block1_addr)));
   LUT_gen23_block2_addr <= allbits(17 downto 12);
   LUT_gen23(2) <= LUT_gen23_block2_data(to_integer(unsigned(LUT_gen23_block2_addr)));
   LUT_gen23_block3_addr <= allbits(23 downto 18);
   LUT_gen23(3) <= LUT_gen23_block3_data(to_integer(unsigned(LUT_gen23_block3_addr)));
   LUT_gen23_block4_addr <= allbits(29 downto 24);
   LUT_gen23(4) <= LUT_gen23_block4_data(to_integer(unsigned(LUT_gen23_block4_addr)));
   LUT_gen23_block5_addr <= allbits(35 downto 30);
   LUT_gen23(5) <= LUT_gen23_block5_data(to_integer(unsigned(LUT_gen23_block5_addr)));
   LUT_gen23_block6_addr <= allbits(41 downto 36);
   LUT_gen23(6) <= LUT_gen23_block6_data(to_integer(unsigned(LUT_gen23_block6_addr)));
   LUT_gen23_block7_addr <= allbits(47 downto 42);
   LUT_gen23(7) <= LUT_gen23_block7_data(to_integer(unsigned(LUT_gen23_block7_addr)));
   LUT_gen23_block8_addr <= allbits(53 downto 48);
   LUT_gen23(8) <= LUT_gen23_block8_data(to_integer(unsigned(LUT_gen23_block8_addr)));
   LUT_gen23_block9_addr <= allbits(59 downto 54);
   LUT_gen23(9) <= LUT_gen23_block9_data(to_integer(unsigned(LUT_gen23_block9_addr)));
   LUT_gen23_block10_addr <= allbits(65 downto 60);
   LUT_gen23(10) <= LUT_gen23_block10_data(to_integer(unsigned(LUT_gen23_block10_addr)));
   LUT_gen23_block11_addr <= allbits(71 downto 66);
   LUT_gen23(11) <= LUT_gen23_block11_data(to_integer(unsigned(LUT_gen23_block11_addr)));
   LUT_gen23_block12_addr <= allbits(77 downto 72);
   LUT_gen23(12) <= LUT_gen23_block12_data(to_integer(unsigned(LUT_gen23_block12_addr)));
   LUT_gen23_block13_addr <= allbits(83 downto 78);
   LUT_gen23(13) <= LUT_gen23_block13_data(to_integer(unsigned(LUT_gen23_block13_addr)));
   LUT_gen23_block14_addr <= allbits(89 downto 84);
   LUT_gen23(14) <= LUT_gen23_block14_data(to_integer(unsigned(LUT_gen23_block14_addr)));
   LUT_gen23_block15_addr <= allbits(95 downto 90);
   LUT_gen23(15) <= LUT_gen23_block15_data(to_integer(unsigned(LUT_gen23_block15_addr)));
   LUT_gen24_block0_addr <= allbits(5 downto 0);
   LUT_gen24(0) <= LUT_gen24_block0_data(to_integer(unsigned(LUT_gen24_block0_addr)));
   LUT_gen24_block1_addr <= allbits(11 downto 6);
   LUT_gen24(1) <= LUT_gen24_block1_data(to_integer(unsigned(LUT_gen24_block1_addr)));
   LUT_gen24_block2_addr <= allbits(17 downto 12);
   LUT_gen24(2) <= LUT_gen24_block2_data(to_integer(unsigned(LUT_gen24_block2_addr)));
   LUT_gen24_block3_addr <= allbits(23 downto 18);
   LUT_gen24(3) <= LUT_gen24_block3_data(to_integer(unsigned(LUT_gen24_block3_addr)));
   LUT_gen24_block4_addr <= allbits(29 downto 24);
   LUT_gen24(4) <= LUT_gen24_block4_data(to_integer(unsigned(LUT_gen24_block4_addr)));
   LUT_gen24_block5_addr <= allbits(35 downto 30);
   LUT_gen24(5) <= LUT_gen24_block5_data(to_integer(unsigned(LUT_gen24_block5_addr)));
   LUT_gen24_block6_addr <= allbits(41 downto 36);
   LUT_gen24(6) <= LUT_gen24_block6_data(to_integer(unsigned(LUT_gen24_block6_addr)));
   LUT_gen24_block7_addr <= allbits(47 downto 42);
   LUT_gen24(7) <= LUT_gen24_block7_data(to_integer(unsigned(LUT_gen24_block7_addr)));
   LUT_gen24_block8_addr <= allbits(53 downto 48);
   LUT_gen24(8) <= LUT_gen24_block8_data(to_integer(unsigned(LUT_gen24_block8_addr)));
   LUT_gen24_block9_addr <= allbits(59 downto 54);
   LUT_gen24(9) <= LUT_gen24_block9_data(to_integer(unsigned(LUT_gen24_block9_addr)));
   LUT_gen24_block10_addr <= allbits(65 downto 60);
   LUT_gen24(10) <= LUT_gen24_block10_data(to_integer(unsigned(LUT_gen24_block10_addr)));
   LUT_gen24_block11_addr <= allbits(71 downto 66);
   LUT_gen24(11) <= LUT_gen24_block11_data(to_integer(unsigned(LUT_gen24_block11_addr)));
   LUT_gen24_block12_addr <= allbits(77 downto 72);
   LUT_gen24(12) <= LUT_gen24_block12_data(to_integer(unsigned(LUT_gen24_block12_addr)));
   LUT_gen24_block13_addr <= allbits(83 downto 78);
   LUT_gen24(13) <= LUT_gen24_block13_data(to_integer(unsigned(LUT_gen24_block13_addr)));
   LUT_gen24_block14_addr <= allbits(89 downto 84);
   LUT_gen24(14) <= LUT_gen24_block14_data(to_integer(unsigned(LUT_gen24_block14_addr)));
   LUT_gen24_block15_addr <= allbits(95 downto 90);
   LUT_gen24(15) <= LUT_gen24_block15_data(to_integer(unsigned(LUT_gen24_block15_addr)));
   LUT_gen25_block0_addr <= allbits(5 downto 0);
   LUT_gen25(0) <= LUT_gen25_block0_data(to_integer(unsigned(LUT_gen25_block0_addr)));
   LUT_gen25_block1_addr <= allbits(11 downto 6);
   LUT_gen25(1) <= LUT_gen25_block1_data(to_integer(unsigned(LUT_gen25_block1_addr)));
   LUT_gen25_block2_addr <= allbits(17 downto 12);
   LUT_gen25(2) <= LUT_gen25_block2_data(to_integer(unsigned(LUT_gen25_block2_addr)));
   LUT_gen25_block3_addr <= allbits(23 downto 18);
   LUT_gen25(3) <= LUT_gen25_block3_data(to_integer(unsigned(LUT_gen25_block3_addr)));
   LUT_gen25_block4_addr <= allbits(29 downto 24);
   LUT_gen25(4) <= LUT_gen25_block4_data(to_integer(unsigned(LUT_gen25_block4_addr)));
   LUT_gen25_block5_addr <= allbits(35 downto 30);
   LUT_gen25(5) <= LUT_gen25_block5_data(to_integer(unsigned(LUT_gen25_block5_addr)));
   LUT_gen25_block6_addr <= allbits(41 downto 36);
   LUT_gen25(6) <= LUT_gen25_block6_data(to_integer(unsigned(LUT_gen25_block6_addr)));
   LUT_gen25_block7_addr <= allbits(47 downto 42);
   LUT_gen25(7) <= LUT_gen25_block7_data(to_integer(unsigned(LUT_gen25_block7_addr)));
   LUT_gen25_block8_addr <= allbits(53 downto 48);
   LUT_gen25(8) <= LUT_gen25_block8_data(to_integer(unsigned(LUT_gen25_block8_addr)));
   LUT_gen25_block9_addr <= allbits(59 downto 54);
   LUT_gen25(9) <= LUT_gen25_block9_data(to_integer(unsigned(LUT_gen25_block9_addr)));
   LUT_gen25_block10_addr <= allbits(65 downto 60);
   LUT_gen25(10) <= LUT_gen25_block10_data(to_integer(unsigned(LUT_gen25_block10_addr)));
   LUT_gen25_block11_addr <= allbits(71 downto 66);
   LUT_gen25(11) <= LUT_gen25_block11_data(to_integer(unsigned(LUT_gen25_block11_addr)));
   LUT_gen25_block12_addr <= allbits(77 downto 72);
   LUT_gen25(12) <= LUT_gen25_block12_data(to_integer(unsigned(LUT_gen25_block12_addr)));
   LUT_gen25_block13_addr <= allbits(83 downto 78);
   LUT_gen25(13) <= LUT_gen25_block13_data(to_integer(unsigned(LUT_gen25_block13_addr)));
   LUT_gen25_block14_addr <= allbits(89 downto 84);
   LUT_gen25(14) <= LUT_gen25_block14_data(to_integer(unsigned(LUT_gen25_block14_addr)));
   LUT_gen25_block15_addr <= allbits(95 downto 90);
   LUT_gen25(15) <= LUT_gen25_block15_data(to_integer(unsigned(LUT_gen25_block15_addr)));
   LUT_gen26_block0_addr <= allbits(5 downto 0);
   LUT_gen26(0) <= LUT_gen26_block0_data(to_integer(unsigned(LUT_gen26_block0_addr)));
   LUT_gen26_block1_addr <= allbits(11 downto 6);
   LUT_gen26(1) <= LUT_gen26_block1_data(to_integer(unsigned(LUT_gen26_block1_addr)));
   LUT_gen26_block2_addr <= allbits(17 downto 12);
   LUT_gen26(2) <= LUT_gen26_block2_data(to_integer(unsigned(LUT_gen26_block2_addr)));
   LUT_gen26_block3_addr <= allbits(23 downto 18);
   LUT_gen26(3) <= LUT_gen26_block3_data(to_integer(unsigned(LUT_gen26_block3_addr)));
   LUT_gen26_block4_addr <= allbits(29 downto 24);
   LUT_gen26(4) <= LUT_gen26_block4_data(to_integer(unsigned(LUT_gen26_block4_addr)));
   LUT_gen26_block5_addr <= allbits(35 downto 30);
   LUT_gen26(5) <= LUT_gen26_block5_data(to_integer(unsigned(LUT_gen26_block5_addr)));
   LUT_gen26_block6_addr <= allbits(41 downto 36);
   LUT_gen26(6) <= LUT_gen26_block6_data(to_integer(unsigned(LUT_gen26_block6_addr)));
   LUT_gen26_block7_addr <= allbits(47 downto 42);
   LUT_gen26(7) <= LUT_gen26_block7_data(to_integer(unsigned(LUT_gen26_block7_addr)));
   LUT_gen26_block8_addr <= allbits(53 downto 48);
   LUT_gen26(8) <= LUT_gen26_block8_data(to_integer(unsigned(LUT_gen26_block8_addr)));
   LUT_gen26_block9_addr <= allbits(59 downto 54);
   LUT_gen26(9) <= LUT_gen26_block9_data(to_integer(unsigned(LUT_gen26_block9_addr)));
   LUT_gen26(10) <= '0';
   LUT_gen26_block11_addr <= allbits(71 downto 66);
   LUT_gen26(11) <= LUT_gen26_block11_data(to_integer(unsigned(LUT_gen26_block11_addr)));
   LUT_gen26_block12_addr <= allbits(77 downto 72);
   LUT_gen26(12) <= LUT_gen26_block12_data(to_integer(unsigned(LUT_gen26_block12_addr)));
   LUT_gen26_block13_addr <= allbits(83 downto 78);
   LUT_gen26(13) <= LUT_gen26_block13_data(to_integer(unsigned(LUT_gen26_block13_addr)));
   LUT_gen26_block14_addr <= allbits(89 downto 84);
   LUT_gen26(14) <= LUT_gen26_block14_data(to_integer(unsigned(LUT_gen26_block14_addr)));
   LUT_gen26_block15_addr <= allbits(95 downto 90);
   LUT_gen26(15) <= LUT_gen26_block15_data(to_integer(unsigned(LUT_gen26_block15_addr)));
   LUT_gen27_block0_addr <= allbits(5 downto 0);
   LUT_gen27(0) <= LUT_gen27_block0_data(to_integer(unsigned(LUT_gen27_block0_addr)));
   LUT_gen27_block1_addr <= allbits(11 downto 6);
   LUT_gen27(1) <= LUT_gen27_block1_data(to_integer(unsigned(LUT_gen27_block1_addr)));
   LUT_gen27_block2_addr <= allbits(17 downto 12);
   LUT_gen27(2) <= LUT_gen27_block2_data(to_integer(unsigned(LUT_gen27_block2_addr)));
   LUT_gen27_block3_addr <= allbits(23 downto 18);
   LUT_gen27(3) <= LUT_gen27_block3_data(to_integer(unsigned(LUT_gen27_block3_addr)));
   LUT_gen27_block4_addr <= allbits(29 downto 24);
   LUT_gen27(4) <= LUT_gen27_block4_data(to_integer(unsigned(LUT_gen27_block4_addr)));
   LUT_gen27_block5_addr <= allbits(35 downto 30);
   LUT_gen27(5) <= LUT_gen27_block5_data(to_integer(unsigned(LUT_gen27_block5_addr)));
   LUT_gen27_block6_addr <= allbits(41 downto 36);
   LUT_gen27(6) <= LUT_gen27_block6_data(to_integer(unsigned(LUT_gen27_block6_addr)));
   LUT_gen27_block7_addr <= allbits(47 downto 42);
   LUT_gen27(7) <= LUT_gen27_block7_data(to_integer(unsigned(LUT_gen27_block7_addr)));
   LUT_gen27_block8_addr <= allbits(53 downto 48);
   LUT_gen27(8) <= LUT_gen27_block8_data(to_integer(unsigned(LUT_gen27_block8_addr)));
   LUT_gen27_block9_addr <= allbits(59 downto 54);
   LUT_gen27(9) <= LUT_gen27_block9_data(to_integer(unsigned(LUT_gen27_block9_addr)));
   LUT_gen27_block10_addr <= allbits(65 downto 60);
   LUT_gen27(10) <= LUT_gen27_block10_data(to_integer(unsigned(LUT_gen27_block10_addr)));
   LUT_gen27_block11_addr <= allbits(71 downto 66);
   LUT_gen27(11) <= LUT_gen27_block11_data(to_integer(unsigned(LUT_gen27_block11_addr)));
   LUT_gen27_block12_addr <= allbits(77 downto 72);
   LUT_gen27(12) <= LUT_gen27_block12_data(to_integer(unsigned(LUT_gen27_block12_addr)));
   LUT_gen27_block13_addr <= allbits(83 downto 78);
   LUT_gen27(13) <= LUT_gen27_block13_data(to_integer(unsigned(LUT_gen27_block13_addr)));
   LUT_gen27_block14_addr <= allbits(89 downto 84);
   LUT_gen27(14) <= LUT_gen27_block14_data(to_integer(unsigned(LUT_gen27_block14_addr)));
   LUT_gen27_block15_addr <= allbits(95 downto 90);
   LUT_gen27(15) <= LUT_gen27_block15_data(to_integer(unsigned(LUT_gen27_block15_addr)));
   LUT_gen28_block0_addr <= allbits(5 downto 0);
   LUT_gen28(0) <= LUT_gen28_block0_data(to_integer(unsigned(LUT_gen28_block0_addr)));
   LUT_gen28_block1_addr <= allbits(11 downto 6);
   LUT_gen28(1) <= LUT_gen28_block1_data(to_integer(unsigned(LUT_gen28_block1_addr)));
   LUT_gen28(2) <= '0';
   LUT_gen28_block3_addr <= allbits(23 downto 18);
   LUT_gen28(3) <= LUT_gen28_block3_data(to_integer(unsigned(LUT_gen28_block3_addr)));
   LUT_gen28_block4_addr <= allbits(29 downto 24);
   LUT_gen28(4) <= LUT_gen28_block4_data(to_integer(unsigned(LUT_gen28_block4_addr)));
   LUT_gen28_block5_addr <= allbits(35 downto 30);
   LUT_gen28(5) <= LUT_gen28_block5_data(to_integer(unsigned(LUT_gen28_block5_addr)));
   LUT_gen28_block6_addr <= allbits(41 downto 36);
   LUT_gen28(6) <= LUT_gen28_block6_data(to_integer(unsigned(LUT_gen28_block6_addr)));
   LUT_gen28_block7_addr <= allbits(47 downto 42);
   LUT_gen28(7) <= LUT_gen28_block7_data(to_integer(unsigned(LUT_gen28_block7_addr)));
   LUT_gen28_block8_addr <= allbits(53 downto 48);
   LUT_gen28(8) <= LUT_gen28_block8_data(to_integer(unsigned(LUT_gen28_block8_addr)));
   LUT_gen28_block9_addr <= allbits(59 downto 54);
   LUT_gen28(9) <= LUT_gen28_block9_data(to_integer(unsigned(LUT_gen28_block9_addr)));
   LUT_gen28_block10_addr <= allbits(65 downto 60);
   LUT_gen28(10) <= LUT_gen28_block10_data(to_integer(unsigned(LUT_gen28_block10_addr)));
   LUT_gen28_block11_addr <= allbits(71 downto 66);
   LUT_gen28(11) <= LUT_gen28_block11_data(to_integer(unsigned(LUT_gen28_block11_addr)));
   LUT_gen28_block12_addr <= allbits(77 downto 72);
   LUT_gen28(12) <= LUT_gen28_block12_data(to_integer(unsigned(LUT_gen28_block12_addr)));
   LUT_gen28_block13_addr <= allbits(83 downto 78);
   LUT_gen28(13) <= LUT_gen28_block13_data(to_integer(unsigned(LUT_gen28_block13_addr)));
   LUT_gen28_block14_addr <= allbits(89 downto 84);
   LUT_gen28(14) <= LUT_gen28_block14_data(to_integer(unsigned(LUT_gen28_block14_addr)));
   LUT_gen28_block15_addr <= allbits(95 downto 90);
   LUT_gen28(15) <= LUT_gen28_block15_data(to_integer(unsigned(LUT_gen28_block15_addr)));
   LUT_gen29_block0_addr <= allbits(5 downto 0);
   LUT_gen29(0) <= LUT_gen29_block0_data(to_integer(unsigned(LUT_gen29_block0_addr)));
   LUT_gen29_block1_addr <= allbits(11 downto 6);
   LUT_gen29(1) <= LUT_gen29_block1_data(to_integer(unsigned(LUT_gen29_block1_addr)));
   LUT_gen29_block2_addr <= allbits(17 downto 12);
   LUT_gen29(2) <= LUT_gen29_block2_data(to_integer(unsigned(LUT_gen29_block2_addr)));
   LUT_gen29_block3_addr <= allbits(23 downto 18);
   LUT_gen29(3) <= LUT_gen29_block3_data(to_integer(unsigned(LUT_gen29_block3_addr)));
   LUT_gen29_block4_addr <= allbits(29 downto 24);
   LUT_gen29(4) <= LUT_gen29_block4_data(to_integer(unsigned(LUT_gen29_block4_addr)));
   LUT_gen29_block5_addr <= allbits(35 downto 30);
   LUT_gen29(5) <= LUT_gen29_block5_data(to_integer(unsigned(LUT_gen29_block5_addr)));
   LUT_gen29_block6_addr <= allbits(41 downto 36);
   LUT_gen29(6) <= LUT_gen29_block6_data(to_integer(unsigned(LUT_gen29_block6_addr)));
   LUT_gen29_block7_addr <= allbits(47 downto 42);
   LUT_gen29(7) <= LUT_gen29_block7_data(to_integer(unsigned(LUT_gen29_block7_addr)));
   LUT_gen29_block8_addr <= allbits(53 downto 48);
   LUT_gen29(8) <= LUT_gen29_block8_data(to_integer(unsigned(LUT_gen29_block8_addr)));
   LUT_gen29_block9_addr <= allbits(59 downto 54);
   LUT_gen29(9) <= LUT_gen29_block9_data(to_integer(unsigned(LUT_gen29_block9_addr)));
   LUT_gen29_block10_addr <= allbits(65 downto 60);
   LUT_gen29(10) <= LUT_gen29_block10_data(to_integer(unsigned(LUT_gen29_block10_addr)));
   LUT_gen29_block11_addr <= allbits(71 downto 66);
   LUT_gen29(11) <= LUT_gen29_block11_data(to_integer(unsigned(LUT_gen29_block11_addr)));
   LUT_gen29_block12_addr <= allbits(77 downto 72);
   LUT_gen29(12) <= LUT_gen29_block12_data(to_integer(unsigned(LUT_gen29_block12_addr)));
   LUT_gen29_block13_addr <= allbits(83 downto 78);
   LUT_gen29(13) <= LUT_gen29_block13_data(to_integer(unsigned(LUT_gen29_block13_addr)));
   LUT_gen29_block14_addr <= allbits(89 downto 84);
   LUT_gen29(14) <= LUT_gen29_block14_data(to_integer(unsigned(LUT_gen29_block14_addr)));
   LUT_gen29_block15_addr <= allbits(95 downto 90);
   LUT_gen29(15) <= LUT_gen29_block15_data(to_integer(unsigned(LUT_gen29_block15_addr)));
   LUT_gen30_block0_addr <= allbits(5 downto 0);
   LUT_gen30(0) <= LUT_gen30_block0_data(to_integer(unsigned(LUT_gen30_block0_addr)));
   LUT_gen30_block1_addr <= allbits(11 downto 6);
   LUT_gen30(1) <= LUT_gen30_block1_data(to_integer(unsigned(LUT_gen30_block1_addr)));
   LUT_gen30_block2_addr <= allbits(17 downto 12);
   LUT_gen30(2) <= LUT_gen30_block2_data(to_integer(unsigned(LUT_gen30_block2_addr)));
   LUT_gen30_block3_addr <= allbits(23 downto 18);
   LUT_gen30(3) <= LUT_gen30_block3_data(to_integer(unsigned(LUT_gen30_block3_addr)));
   LUT_gen30_block4_addr <= allbits(29 downto 24);
   LUT_gen30(4) <= LUT_gen30_block4_data(to_integer(unsigned(LUT_gen30_block4_addr)));
   LUT_gen30_block5_addr <= allbits(35 downto 30);
   LUT_gen30(5) <= LUT_gen30_block5_data(to_integer(unsigned(LUT_gen30_block5_addr)));
   LUT_gen30_block6_addr <= allbits(41 downto 36);
   LUT_gen30(6) <= LUT_gen30_block6_data(to_integer(unsigned(LUT_gen30_block6_addr)));
   LUT_gen30_block7_addr <= allbits(47 downto 42);
   LUT_gen30(7) <= LUT_gen30_block7_data(to_integer(unsigned(LUT_gen30_block7_addr)));
   LUT_gen30_block8_addr <= allbits(53 downto 48);
   LUT_gen30(8) <= LUT_gen30_block8_data(to_integer(unsigned(LUT_gen30_block8_addr)));
   LUT_gen30_block9_addr <= allbits(59 downto 54);
   LUT_gen30(9) <= LUT_gen30_block9_data(to_integer(unsigned(LUT_gen30_block9_addr)));
   LUT_gen30_block10_addr <= allbits(65 downto 60);
   LUT_gen30(10) <= LUT_gen30_block10_data(to_integer(unsigned(LUT_gen30_block10_addr)));
   LUT_gen30_block11_addr <= allbits(71 downto 66);
   LUT_gen30(11) <= LUT_gen30_block11_data(to_integer(unsigned(LUT_gen30_block11_addr)));
   LUT_gen30(12) <= '0';
   LUT_gen30_block13_addr <= allbits(83 downto 78);
   LUT_gen30(13) <= LUT_gen30_block13_data(to_integer(unsigned(LUT_gen30_block13_addr)));
   LUT_gen30_block14_addr <= allbits(89 downto 84);
   LUT_gen30(14) <= LUT_gen30_block14_data(to_integer(unsigned(LUT_gen30_block14_addr)));
   LUT_gen30_block15_addr <= allbits(95 downto 90);
   LUT_gen30(15) <= LUT_gen30_block15_data(to_integer(unsigned(LUT_gen30_block15_addr)));
   LUT_gen31_block0_addr <= allbits(5 downto 0);
   LUT_gen31(0) <= LUT_gen31_block0_data(to_integer(unsigned(LUT_gen31_block0_addr)));
   LUT_gen31_block1_addr <= allbits(11 downto 6);
   LUT_gen31(1) <= LUT_gen31_block1_data(to_integer(unsigned(LUT_gen31_block1_addr)));
   LUT_gen31_block2_addr <= allbits(17 downto 12);
   LUT_gen31(2) <= LUT_gen31_block2_data(to_integer(unsigned(LUT_gen31_block2_addr)));
   LUT_gen31_block3_addr <= allbits(23 downto 18);
   LUT_gen31(3) <= LUT_gen31_block3_data(to_integer(unsigned(LUT_gen31_block3_addr)));
   LUT_gen31_block4_addr <= allbits(29 downto 24);
   LUT_gen31(4) <= LUT_gen31_block4_data(to_integer(unsigned(LUT_gen31_block4_addr)));
   LUT_gen31_block5_addr <= allbits(35 downto 30);
   LUT_gen31(5) <= LUT_gen31_block5_data(to_integer(unsigned(LUT_gen31_block5_addr)));
   LUT_gen31_block6_addr <= allbits(41 downto 36);
   LUT_gen31(6) <= LUT_gen31_block6_data(to_integer(unsigned(LUT_gen31_block6_addr)));
   LUT_gen31_block7_addr <= allbits(47 downto 42);
   LUT_gen31(7) <= LUT_gen31_block7_data(to_integer(unsigned(LUT_gen31_block7_addr)));
   LUT_gen31_block8_addr <= allbits(53 downto 48);
   LUT_gen31(8) <= LUT_gen31_block8_data(to_integer(unsigned(LUT_gen31_block8_addr)));
   LUT_gen31_block9_addr <= allbits(59 downto 54);
   LUT_gen31(9) <= LUT_gen31_block9_data(to_integer(unsigned(LUT_gen31_block9_addr)));
   LUT_gen31_block10_addr <= allbits(65 downto 60);
   LUT_gen31(10) <= LUT_gen31_block10_data(to_integer(unsigned(LUT_gen31_block10_addr)));
   LUT_gen31_block11_addr <= allbits(71 downto 66);
   LUT_gen31(11) <= LUT_gen31_block11_data(to_integer(unsigned(LUT_gen31_block11_addr)));
   LUT_gen31(12) <= '0';
   LUT_gen31_block13_addr <= allbits(83 downto 78);
   LUT_gen31(13) <= LUT_gen31_block13_data(to_integer(unsigned(LUT_gen31_block13_addr)));
   LUT_gen31_block14_addr <= allbits(89 downto 84);
   LUT_gen31(14) <= LUT_gen31_block14_data(to_integer(unsigned(LUT_gen31_block14_addr)));
   LUT_gen31_block15_addr <= allbits(95 downto 90);
   LUT_gen31(15) <= LUT_gen31_block15_data(to_integer(unsigned(LUT_gen31_block15_addr)));

end Behavioral;
