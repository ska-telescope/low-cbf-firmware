LIBRARY IEEE, technology_lib;
USE IEEE.std_logic_1164.ALL;
USE technology_lib.technology_pkg.ALL;


PACKAGE tech_hbm_pkg IS

   TYPE t_hbm_configuration IS (
      HBM_CONFIG_LEFT_FULL, HBM_CONFIG_RIGHT_INDIVIDUAL);




END tech_hbm_pkg;

