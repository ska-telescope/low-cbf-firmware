--------------------------------------------------------------------------------
-- Copyright (C) 1999-2008 Easics NV.
-- This source file may be used and distributed without restriction
-- provided that this copyright statement is not removed from the file
-- and that any derivative work contains the original copyright notice
-- and the associated disclaimer.
--
-- THIS SOURCE FILE IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS
-- OR IMPLIED WARRANTIES, INCLUDING, WITHOUT LIMITATION, THE IMPLIED
-- WARRANTIES OF MERCHANTIBILITY AND FITNESS FOR A PARTICULAR PURPOSE.
--
-- Purpose : synthesizable CRC function
--   * polynomial: (0 1 2 4 5 7 8 10 11 12 16 22 23 26 32)
--   * data width: 512
--
-- Info : tools@easics.be
--        http://www.easics.com
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

package PCK_CRC32_D512 is
  -- polynomial: (0 1 2 4 5 7 8 10 11 12 16 22 23 26 32)
  -- data width: 512
  -- convention: the first serial bit is D[511]
  function nextCRC32_D512
    (Data: std_logic_vector(511 downto 0);
     crc:  std_logic_vector(31 downto 0))
    return std_logic_vector;
end PCK_CRC32_D512;


package body PCK_CRC32_D512 is

  -- polynomial: (0 1 2 4 5 7 8 10 11 12 16 22 23 26 32)
  -- data width: 512
  -- convention: the first serial bit is D[511]
  function nextCRC32_D512
    (Data: std_logic_vector(511 downto 0);
     crc:  std_logic_vector(31 downto 0))
    return std_logic_vector is

    variable d:      std_logic_vector(511 downto 0);
    variable c:      std_logic_vector(31 downto 0);
    variable newcrc: std_logic_vector(31 downto 0);

  begin
    d := Data;
    c := crc;

    newcrc(0) := d(511) xor d(510) xor d(508) xor d(507) xor d(506) xor d(502) xor d(501) xor d(500) xor d(495) xor d(494) xor d(493) xor d(492) xor d(491) xor d(490) xor d(489) xor d(488) xor d(486) xor d(483) xor d(482) xor d(481) xor d(480) xor d(479) xor d(477) xor d(476) xor d(472) xor d(470) xor d(468) xor d(465) xor d(464) xor d(462) xor d(461) xor d(458) xor d(452) xor d(450) xor d(449) xor d(448) xor d(444) xor d(437) xor d(436) xor d(434) xor d(433) xor d(424) xor d(422) xor d(419) xor d(418) xor d(416) xor d(414) xor d(412) xor d(409) xor d(408) xor d(407) xor d(405) xor d(404) xor d(400) xor d(399) xor d(398) xor d(396) xor d(393) xor d(392) xor d(391) xor d(390) xor d(388) xor d(387) xor d(386) xor d(381) xor d(378) xor d(376) xor d(374) xor d(372) xor d(369) xor d(368) xor d(366) xor d(363) xor d(362) xor d(359) xor d(358) xor d(357) xor d(353) xor d(349) xor d(348) xor d(347) xor d(345) xor d(344) xor d(342) xor d(341) xor d(339) xor d(338) xor d(337) xor d(335) xor d(334) xor d(333) xor d(328) xor d(327) xor d(322) xor d(321) xor d(320) xor d(319) xor d(318) xor d(317) xor d(315) xor d(312) xor d(310) xor d(309) xor d(305) xor d(303) xor d(302) xor d(300) xor d(299) xor d(298) xor d(297) xor d(296) xor d(295) xor d(294) xor d(292) xor d(290) xor d(288) xor d(287) xor d(286) xor d(283) xor d(279) xor d(277) xor d(276) xor d(274) xor d(273) xor d(269) xor d(268) xor d(265) xor d(264) xor d(261) xor d(259) xor d(257) xor d(255) xor d(252) xor d(248) xor d(243) xor d(237) xor d(234) xor d(230) xor d(228) xor d(227) xor d(226) xor d(224) xor d(216) xor d(214) xor d(212) xor d(210) xor d(209) xor d(208) xor d(207) xor d(203) xor d(202) xor d(201) xor d(199) xor d(198) xor d(197) xor d(194) xor d(193) xor d(192) xor d(191) xor d(190) xor d(188) xor d(186) xor d(183) xor d(182) xor d(172) xor d(171) xor d(170) xor d(169) xor d(167) xor d(166) xor d(162) xor d(161) xor d(158) xor d(156) xor d(155) xor d(151) xor d(149) xor d(144) xor d(143) xor d(137) xor d(136) xor d(135) xor d(134) xor d(132) xor d(128) xor d(127) xor d(126) xor d(125) xor d(123) xor d(119) xor d(118) xor d(117) xor d(116) xor d(114) xor d(113) xor d(111) xor d(110) xor d(106) xor d(104) xor d(103) xor d(101) xor d(99) xor d(98) xor d(97) xor d(96) xor d(95) xor d(94) xor d(87) xor d(85) xor d(84) xor d(83) xor d(82) xor d(81) xor d(79) xor d(73) xor d(72) xor d(68) xor d(67) xor d(66) xor d(65) xor d(63) xor d(61) xor d(60) xor d(58) xor d(55) xor d(54) xor d(53) xor d(50) xor d(48) xor d(47) xor d(45) xor d(44) xor d(37) xor d(34) xor d(32) xor d(31) xor d(30) xor d(29) xor d(28) xor d(26) xor d(25) xor d(24) xor d(16) xor d(12) xor d(10) xor d(9) xor d(6) xor d(0) xor c(0) xor c(1) xor c(2) xor c(3) xor c(6) xor c(8) xor c(9) xor c(10) xor c(11) xor c(12) xor c(13) xor c(14) xor c(15) xor c(20) xor c(21) xor c(22) xor c(26) xor c(27) xor c(28) xor c(30) xor c(31);
    newcrc(1) := d(510) xor d(509) xor d(506) xor d(503) xor d(500) xor d(496) xor d(488) xor d(487) xor d(486) xor d(484) xor d(479) xor d(478) xor d(476) xor d(473) xor d(472) xor d(471) xor d(470) xor d(469) xor d(468) xor d(466) xor d(464) xor d(463) xor d(461) xor d(459) xor d(458) xor d(453) xor d(452) xor d(451) xor d(448) xor d(445) xor d(444) xor d(438) xor d(436) xor d(435) xor d(433) xor d(425) xor d(424) xor d(423) xor d(422) xor d(420) xor d(418) xor d(417) xor d(416) xor d(415) xor d(414) xor d(413) xor d(412) xor d(410) xor d(407) xor d(406) xor d(404) xor d(401) xor d(398) xor d(397) xor d(396) xor d(394) xor d(390) xor d(389) xor d(386) xor d(382) xor d(381) xor d(379) xor d(378) xor d(377) xor d(376) xor d(375) xor d(374) xor d(373) xor d(372) xor d(370) xor d(368) xor d(367) xor d(366) xor d(364) xor d(362) xor d(360) xor d(357) xor d(354) xor d(353) xor d(350) xor d(347) xor d(346) xor d(344) xor d(343) xor d(341) xor d(340) xor d(337) xor d(336) xor d(333) xor d(329) xor d(327) xor d(323) xor d(317) xor d(316) xor d(315) xor d(313) xor d(312) xor d(311) xor d(309) xor d(306) xor d(305) xor d(304) xor d(302) xor d(301) xor d(294) xor d(293) xor d(292) xor d(291) xor d(290) xor d(289) xor d(286) xor d(284) xor d(283) xor d(280) xor d(279) xor d(278) xor d(276) xor d(275) xor d(273) xor d(270) xor d(268) xor d(266) xor d(264) xor d(262) xor d(261) xor d(260) xor d(259) xor d(258) xor d(257) xor d(256) xor d(255) xor d(253) xor d(252) xor d(249) xor d(248) xor d(244) xor d(243) xor d(238) xor d(237) xor d(235) xor d(234) xor d(231) xor d(230) xor d(229) xor d(226) xor d(225) xor d(224) xor d(217) xor d(216) xor d(215) xor d(214) xor d(213) xor d(212) xor d(211) xor d(207) xor d(204) xor d(201) xor d(200) xor d(197) xor d(195) xor d(190) xor d(189) xor d(188) xor d(187) xor d(186) xor d(184) xor d(182) xor d(173) xor d(169) xor d(168) xor d(166) xor d(163) xor d(161) xor d(159) xor d(158) xor d(157) xor d(155) xor d(152) xor d(151) xor d(150) xor d(149) xor d(145) xor d(143) xor d(138) xor d(134) xor d(133) xor d(132) xor d(129) xor d(125) xor d(124) xor d(123) xor d(120) xor d(116) xor d(115) xor d(113) xor d(112) xor d(110) xor d(107) xor d(106) xor d(105) xor d(103) xor d(102) xor d(101) xor d(100) xor d(94) xor d(88) xor d(87) xor d(86) xor d(81) xor d(80) xor d(79) xor d(74) xor d(72) xor d(69) xor d(65) xor d(64) xor d(63) xor d(62) xor d(60) xor d(59) xor d(58) xor d(56) xor d(53) xor d(51) xor d(50) xor d(49) xor d(47) xor d(46) xor d(44) xor d(38) xor d(37) xor d(35) xor d(34) xor d(33) xor d(28) xor d(27) xor d(24) xor d(17) xor d(16) xor d(13) xor d(12) xor d(11) xor d(9) xor d(7) xor d(6) xor d(1) xor d(0) xor c(4) xor c(6) xor c(7) xor c(8) xor c(16) xor c(20) xor c(23) xor c(26) xor c(29) xor c(30);
    newcrc(2) := d(508) xor d(506) xor d(504) xor d(502) xor d(500) xor d(497) xor d(495) xor d(494) xor d(493) xor d(492) xor d(491) xor d(490) xor d(487) xor d(486) xor d(485) xor d(483) xor d(482) xor d(481) xor d(476) xor d(474) xor d(473) xor d(471) xor d(469) xor d(468) xor d(467) xor d(461) xor d(460) xor d(459) xor d(458) xor d(454) xor d(453) xor d(450) xor d(448) xor d(446) xor d(445) xor d(444) xor d(439) xor d(433) xor d(426) xor d(425) xor d(423) xor d(422) xor d(421) xor d(417) xor d(415) xor d(413) xor d(412) xor d(411) xor d(409) xor d(404) xor d(402) xor d(400) xor d(397) xor d(396) xor d(395) xor d(393) xor d(392) xor d(388) xor d(386) xor d(383) xor d(382) xor d(381) xor d(380) xor d(379) xor d(377) xor d(375) xor d(373) xor d(372) xor d(371) xor d(367) xor d(366) xor d(365) xor d(362) xor d(361) xor d(359) xor d(357) xor d(355) xor d(354) xor d(353) xor d(351) xor d(349) xor d(339) xor d(335) xor d(333) xor d(330) xor d(327) xor d(324) xor d(322) xor d(321) xor d(320) xor d(319) xor d(316) xor d(315) xor d(314) xor d(313) xor d(309) xor d(307) xor d(306) xor d(300) xor d(299) xor d(298) xor d(297) xor d(296) xor d(293) xor d(291) xor d(288) xor d(286) xor d(285) xor d(284) xor d(283) xor d(281) xor d(280) xor d(273) xor d(271) xor d(268) xor d(267) xor d(264) xor d(263) xor d(262) xor d(260) xor d(258) xor d(256) xor d(255) xor d(254) xor d(253) xor d(252) xor d(250) xor d(249) xor d(248) xor d(245) xor d(244) xor d(243) xor d(239) xor d(238) xor d(237) xor d(236) xor d(235) xor d(234) xor d(232) xor d(231) xor d(228) xor d(225) xor d(224) xor d(218) xor d(217) xor d(215) xor d(213) xor d(210) xor d(209) xor d(207) xor d(205) xor d(203) xor d(199) xor d(197) xor d(196) xor d(194) xor d(193) xor d(192) xor d(189) xor d(187) xor d(186) xor d(185) xor d(182) xor d(174) xor d(172) xor d(171) xor d(166) xor d(164) xor d(161) xor d(160) xor d(159) xor d(155) xor d(153) xor d(152) xor d(150) xor d(149) xor d(146) xor d(143) xor d(139) xor d(137) xor d(136) xor d(133) xor d(132) xor d(130) xor d(128) xor d(127) xor d(124) xor d(123) xor d(121) xor d(119) xor d(118) xor d(110) xor d(108) xor d(107) xor d(102) xor d(99) xor d(98) xor d(97) xor d(96) xor d(94) xor d(89) xor d(88) xor d(85) xor d(84) xor d(83) xor d(80) xor d(79) xor d(75) xor d(72) xor d(70) xor d(68) xor d(67) xor d(64) xor d(59) xor d(58) xor d(57) xor d(55) xor d(53) xor d(52) xor d(51) xor d(44) xor d(39) xor d(38) xor d(37) xor d(36) xor d(35) xor d(32) xor d(31) xor d(30) xor d(26) xor d(24) xor d(18) xor d(17) xor d(16) xor d(14) xor d(13) xor d(9) xor d(8) xor d(7) xor d(6) xor d(2) xor d(1) xor d(0) xor c(1) xor c(2) xor c(3) xor c(5) xor c(6) xor c(7) xor c(10) xor c(11) xor c(12) xor c(13) xor c(14) xor c(15) xor c(17) xor c(20) xor c(22) xor c(24) xor c(26) xor c(28);
    newcrc(3) := d(509) xor d(507) xor d(505) xor d(503) xor d(501) xor d(498) xor d(496) xor d(495) xor d(494) xor d(493) xor d(492) xor d(491) xor d(488) xor d(487) xor d(486) xor d(484) xor d(483) xor d(482) xor d(477) xor d(475) xor d(474) xor d(472) xor d(470) xor d(469) xor d(468) xor d(462) xor d(461) xor d(460) xor d(459) xor d(455) xor d(454) xor d(451) xor d(449) xor d(447) xor d(446) xor d(445) xor d(440) xor d(434) xor d(427) xor d(426) xor d(424) xor d(423) xor d(422) xor d(418) xor d(416) xor d(414) xor d(413) xor d(412) xor d(410) xor d(405) xor d(403) xor d(401) xor d(398) xor d(397) xor d(396) xor d(394) xor d(393) xor d(389) xor d(387) xor d(384) xor d(383) xor d(382) xor d(381) xor d(380) xor d(378) xor d(376) xor d(374) xor d(373) xor d(372) xor d(368) xor d(367) xor d(366) xor d(363) xor d(362) xor d(360) xor d(358) xor d(356) xor d(355) xor d(354) xor d(352) xor d(350) xor d(340) xor d(336) xor d(334) xor d(331) xor d(328) xor d(325) xor d(323) xor d(322) xor d(321) xor d(320) xor d(317) xor d(316) xor d(315) xor d(314) xor d(310) xor d(308) xor d(307) xor d(301) xor d(300) xor d(299) xor d(298) xor d(297) xor d(294) xor d(292) xor d(289) xor d(287) xor d(286) xor d(285) xor d(284) xor d(282) xor d(281) xor d(274) xor d(272) xor d(269) xor d(268) xor d(265) xor d(264) xor d(263) xor d(261) xor d(259) xor d(257) xor d(256) xor d(255) xor d(254) xor d(253) xor d(251) xor d(250) xor d(249) xor d(246) xor d(245) xor d(244) xor d(240) xor d(239) xor d(238) xor d(237) xor d(236) xor d(235) xor d(233) xor d(232) xor d(229) xor d(226) xor d(225) xor d(219) xor d(218) xor d(216) xor d(214) xor d(211) xor d(210) xor d(208) xor d(206) xor d(204) xor d(200) xor d(198) xor d(197) xor d(195) xor d(194) xor d(193) xor d(190) xor d(188) xor d(187) xor d(186) xor d(183) xor d(175) xor d(173) xor d(172) xor d(167) xor d(165) xor d(162) xor d(161) xor d(160) xor d(156) xor d(154) xor d(153) xor d(151) xor d(150) xor d(147) xor d(144) xor d(140) xor d(138) xor d(137) xor d(134) xor d(133) xor d(131) xor d(129) xor d(128) xor d(125) xor d(124) xor d(122) xor d(120) xor d(119) xor d(111) xor d(109) xor d(108) xor d(103) xor d(100) xor d(99) xor d(98) xor d(97) xor d(95) xor d(90) xor d(89) xor d(86) xor d(85) xor d(84) xor d(81) xor d(80) xor d(76) xor d(73) xor d(71) xor d(69) xor d(68) xor d(65) xor d(60) xor d(59) xor d(58) xor d(56) xor d(54) xor d(53) xor d(52) xor d(45) xor d(40) xor d(39) xor d(38) xor d(37) xor d(36) xor d(33) xor d(32) xor d(31) xor d(27) xor d(25) xor d(19) xor d(18) xor d(17) xor d(15) xor d(14) xor d(10) xor d(9) xor d(8) xor d(7) xor d(3) xor d(2) xor d(1) xor c(2) xor c(3) xor c(4) xor c(6) xor c(7) xor c(8) xor c(11) xor c(12) xor c(13) xor c(14) xor c(15) xor c(16) xor c(18) xor c(21) xor c(23) xor c(25) xor c(27) xor c(29);
    newcrc(4) := d(511) xor d(507) xor d(504) xor d(501) xor d(500) xor d(499) xor d(497) xor d(496) xor d(491) xor d(490) xor d(487) xor d(486) xor d(485) xor d(484) xor d(482) xor d(481) xor d(480) xor d(479) xor d(478) xor d(477) xor d(475) xor d(473) xor d(472) xor d(471) xor d(469) xor d(468) xor d(465) xor d(464) xor d(463) xor d(460) xor d(458) xor d(456) xor d(455) xor d(449) xor d(447) xor d(446) xor d(444) xor d(441) xor d(437) xor d(436) xor d(435) xor d(434) xor d(433) xor d(428) xor d(427) xor d(425) xor d(423) xor d(422) xor d(418) xor d(417) xor d(416) xor d(415) xor d(413) xor d(412) xor d(411) xor d(409) xor d(408) xor d(407) xor d(406) xor d(405) xor d(402) xor d(400) xor d(397) xor d(396) xor d(395) xor d(394) xor d(393) xor d(392) xor d(391) xor d(387) xor d(386) xor d(385) xor d(384) xor d(383) xor d(382) xor d(379) xor d(378) xor d(377) xor d(376) xor d(375) xor d(373) xor d(372) xor d(367) xor d(366) xor d(364) xor d(362) xor d(361) xor d(358) xor d(356) xor d(355) xor d(351) xor d(349) xor d(348) xor d(347) xor d(345) xor d(344) xor d(342) xor d(339) xor d(338) xor d(334) xor d(333) xor d(332) xor d(329) xor d(328) xor d(327) xor d(326) xor d(324) xor d(323) xor d(320) xor d(319) xor d(316) xor d(312) xor d(311) xor d(310) xor d(308) xor d(305) xor d(303) xor d(301) xor d(297) xor d(296) xor d(294) xor d(293) xor d(292) xor d(285) xor d(282) xor d(279) xor d(277) xor d(276) xor d(275) xor d(274) xor d(270) xor d(268) xor d(266) xor d(262) xor d(261) xor d(260) xor d(259) xor d(258) xor d(256) xor d(254) xor d(251) xor d(250) xor d(248) xor d(247) xor d(246) xor d(245) xor d(243) xor d(241) xor d(240) xor d(239) xor d(238) xor d(236) xor d(233) xor d(228) xor d(224) xor d(220) xor d(219) xor d(217) xor d(216) xor d(215) xor d(214) xor d(211) xor d(210) xor d(208) xor d(205) xor d(203) xor d(202) xor d(197) xor d(196) xor d(195) xor d(193) xor d(192) xor d(190) xor d(189) xor d(187) xor d(186) xor d(184) xor d(183) xor d(182) xor d(176) xor d(174) xor d(173) xor d(172) xor d(171) xor d(170) xor d(169) xor d(168) xor d(167) xor d(163) xor d(158) xor d(157) xor d(156) xor d(154) xor d(152) xor d(149) xor d(148) xor d(145) xor d(144) xor d(143) xor d(141) xor d(139) xor d(138) xor d(137) xor d(136) xor d(130) xor d(129) xor d(128) xor d(127) xor d(121) xor d(120) xor d(119) xor d(118) xor d(117) xor d(116) xor d(114) xor d(113) xor d(112) xor d(111) xor d(109) xor d(106) xor d(103) xor d(100) xor d(97) xor d(95) xor d(94) xor d(91) xor d(90) xor d(86) xor d(84) xor d(83) xor d(79) xor d(77) xor d(74) xor d(73) xor d(70) xor d(69) xor d(68) xor d(67) xor d(65) xor d(63) xor d(59) xor d(58) xor d(57) xor d(50) xor d(48) xor d(47) xor d(46) xor d(45) xor d(44) xor d(41) xor d(40) xor d(39) xor d(38) xor d(33) xor d(31) xor d(30) xor d(29) xor d(25) xor d(24) xor d(20) xor d(19) xor d(18) xor d(15) xor d(12) xor d(11) xor d(8) xor d(6) xor d(4) xor d(3) xor d(2) xor d(0) xor c(0) xor c(1) xor c(2) xor c(4) xor c(5) xor c(6) xor c(7) xor c(10) xor c(11) xor c(16) xor c(17) xor c(19) xor c(20) xor c(21) xor c(24) xor c(27) xor c(31);
    newcrc(5) := d(511) xor d(510) xor d(507) xor d(506) xor d(505) xor d(498) xor d(497) xor d(495) xor d(494) xor d(493) xor d(490) xor d(489) xor d(487) xor d(485) xor d(478) xor d(477) xor d(474) xor d(473) xor d(469) xor d(468) xor d(466) xor d(462) xor d(459) xor d(458) xor d(457) xor d(456) xor d(452) xor d(449) xor d(447) xor d(445) xor d(444) xor d(442) xor d(438) xor d(435) xor d(433) xor d(429) xor d(428) xor d(426) xor d(423) xor d(422) xor d(417) xor d(413) xor d(410) xor d(406) xor d(405) xor d(404) xor d(403) xor d(401) xor d(400) xor d(399) xor d(397) xor d(395) xor d(394) xor d(391) xor d(390) xor d(385) xor d(384) xor d(383) xor d(381) xor d(380) xor d(379) xor d(377) xor d(373) xor d(372) xor d(369) xor d(367) xor d(366) xor d(365) xor d(358) xor d(356) xor d(353) xor d(352) xor d(350) xor d(347) xor d(346) xor d(344) xor d(343) xor d(342) xor d(341) xor d(340) xor d(338) xor d(337) xor d(330) xor d(329) xor d(325) xor d(324) xor d(322) xor d(319) xor d(318) xor d(315) xor d(313) xor d(311) xor d(310) xor d(306) xor d(305) xor d(304) xor d(303) xor d(300) xor d(299) xor d(296) xor d(293) xor d(292) xor d(290) xor d(288) xor d(287) xor d(280) xor d(279) xor d(278) xor d(275) xor d(274) xor d(273) xor d(271) xor d(268) xor d(267) xor d(265) xor d(264) xor d(263) xor d(262) xor d(260) xor d(251) xor d(249) xor d(247) xor d(246) xor d(244) xor d(243) xor d(242) xor d(241) xor d(240) xor d(239) xor d(230) xor d(229) xor d(228) xor d(227) xor d(226) xor d(225) xor d(224) xor d(221) xor d(220) xor d(218) xor d(217) xor d(215) xor d(214) xor d(211) xor d(210) xor d(208) xor d(207) xor d(206) xor d(204) xor d(202) xor d(201) xor d(199) xor d(196) xor d(192) xor d(187) xor d(186) xor d(185) xor d(184) xor d(182) xor d(177) xor d(175) xor d(174) xor d(173) xor d(168) xor d(167) xor d(166) xor d(164) xor d(162) xor d(161) xor d(159) xor d(157) xor d(156) xor d(153) xor d(151) xor d(150) xor d(146) xor d(145) xor d(143) xor d(142) xor d(140) xor d(139) xor d(138) xor d(136) xor d(135) xor d(134) xor d(132) xor d(131) xor d(130) xor d(129) xor d(127) xor d(126) xor d(125) xor d(123) xor d(122) xor d(121) xor d(120) xor d(116) xor d(115) xor d(112) xor d(111) xor d(107) xor d(106) xor d(103) xor d(99) xor d(97) xor d(94) xor d(92) xor d(91) xor d(83) xor d(82) xor d(81) xor d(80) xor d(79) xor d(78) xor d(75) xor d(74) xor d(73) xor d(72) xor d(71) xor d(70) xor d(69) xor d(67) xor d(65) xor d(64) xor d(63) xor d(61) xor d(59) xor d(55) xor d(54) xor d(53) xor d(51) xor d(50) xor d(49) xor d(46) xor d(44) xor d(42) xor d(41) xor d(40) xor d(39) xor d(37) xor d(29) xor d(28) xor d(24) xor d(21) xor d(20) xor d(19) xor d(13) xor d(10) xor d(7) xor d(6) xor d(5) xor d(4) xor d(3) xor d(1) xor d(0) xor c(5) xor c(7) xor c(9) xor c(10) xor c(13) xor c(14) xor c(15) xor c(17) xor c(18) xor c(25) xor c(26) xor c(27) xor c(30) xor c(31);
    newcrc(6) := d(511) xor d(508) xor d(507) xor d(506) xor d(499) xor d(498) xor d(496) xor d(495) xor d(494) xor d(491) xor d(490) xor d(488) xor d(486) xor d(479) xor d(478) xor d(475) xor d(474) xor d(470) xor d(469) xor d(467) xor d(463) xor d(460) xor d(459) xor d(458) xor d(457) xor d(453) xor d(450) xor d(448) xor d(446) xor d(445) xor d(443) xor d(439) xor d(436) xor d(434) xor d(430) xor d(429) xor d(427) xor d(424) xor d(423) xor d(418) xor d(414) xor d(411) xor d(407) xor d(406) xor d(405) xor d(404) xor d(402) xor d(401) xor d(400) xor d(398) xor d(396) xor d(395) xor d(392) xor d(391) xor d(386) xor d(385) xor d(384) xor d(382) xor d(381) xor d(380) xor d(378) xor d(374) xor d(373) xor d(370) xor d(368) xor d(367) xor d(366) xor d(359) xor d(357) xor d(354) xor d(353) xor d(351) xor d(348) xor d(347) xor d(345) xor d(344) xor d(343) xor d(342) xor d(341) xor d(339) xor d(338) xor d(331) xor d(330) xor d(326) xor d(325) xor d(323) xor d(320) xor d(319) xor d(316) xor d(314) xor d(312) xor d(311) xor d(307) xor d(306) xor d(305) xor d(304) xor d(301) xor d(300) xor d(297) xor d(294) xor d(293) xor d(291) xor d(289) xor d(288) xor d(281) xor d(280) xor d(279) xor d(276) xor d(275) xor d(274) xor d(272) xor d(269) xor d(268) xor d(266) xor d(265) xor d(264) xor d(263) xor d(261) xor d(252) xor d(250) xor d(248) xor d(247) xor d(245) xor d(244) xor d(243) xor d(242) xor d(241) xor d(240) xor d(231) xor d(230) xor d(229) xor d(228) xor d(227) xor d(226) xor d(225) xor d(222) xor d(221) xor d(219) xor d(218) xor d(216) xor d(215) xor d(212) xor d(211) xor d(209) xor d(208) xor d(207) xor d(205) xor d(203) xor d(202) xor d(200) xor d(197) xor d(193) xor d(188) xor d(187) xor d(186) xor d(185) xor d(183) xor d(178) xor d(176) xor d(175) xor d(174) xor d(169) xor d(168) xor d(167) xor d(165) xor d(163) xor d(162) xor d(160) xor d(158) xor d(157) xor d(154) xor d(152) xor d(151) xor d(147) xor d(146) xor d(144) xor d(143) xor d(141) xor d(140) xor d(139) xor d(137) xor d(136) xor d(135) xor d(133) xor d(132) xor d(131) xor d(130) xor d(128) xor d(127) xor d(126) xor d(124) xor d(123) xor d(122) xor d(121) xor d(117) xor d(116) xor d(113) xor d(112) xor d(108) xor d(107) xor d(104) xor d(100) xor d(98) xor d(95) xor d(93) xor d(92) xor d(84) xor d(83) xor d(82) xor d(81) xor d(80) xor d(79) xor d(76) xor d(75) xor d(74) xor d(73) xor d(72) xor d(71) xor d(70) xor d(68) xor d(66) xor d(65) xor d(64) xor d(62) xor d(60) xor d(56) xor d(55) xor d(54) xor d(52) xor d(51) xor d(50) xor d(47) xor d(45) xor d(43) xor d(42) xor d(41) xor d(40) xor d(38) xor d(30) xor d(29) xor d(25) xor d(22) xor d(21) xor d(20) xor d(14) xor d(11) xor d(8) xor d(7) xor d(6) xor d(5) xor d(4) xor d(2) xor d(1) xor c(6) xor c(8) xor c(10) xor c(11) xor c(14) xor c(15) xor c(16) xor c(18) xor c(19) xor c(26) xor c(27) xor c(28) xor c(31);
    newcrc(7) := d(511) xor d(510) xor d(509) xor d(506) xor d(502) xor d(501) xor d(499) xor d(497) xor d(496) xor d(494) xor d(493) xor d(490) xor d(488) xor d(487) xor d(486) xor d(483) xor d(482) xor d(481) xor d(477) xor d(475) xor d(472) xor d(471) xor d(465) xor d(462) xor d(460) xor d(459) xor d(454) xor d(452) xor d(451) xor d(450) xor d(448) xor d(447) xor d(446) xor d(440) xor d(436) xor d(435) xor d(434) xor d(433) xor d(431) xor d(430) xor d(428) xor d(425) xor d(422) xor d(418) xor d(416) xor d(415) xor d(414) xor d(409) xor d(406) xor d(404) xor d(403) xor d(402) xor d(401) xor d(400) xor d(398) xor d(397) xor d(391) xor d(390) xor d(388) xor d(385) xor d(383) xor d(382) xor d(379) xor d(378) xor d(376) xor d(375) xor d(372) xor d(371) xor d(367) xor d(366) xor d(363) xor d(362) xor d(360) xor d(359) xor d(357) xor d(355) xor d(354) xor d(353) xor d(352) xor d(347) xor d(346) xor d(343) xor d(341) xor d(340) xor d(338) xor d(337) xor d(335) xor d(334) xor d(333) xor d(332) xor d(331) xor d(328) xor d(326) xor d(324) xor d(322) xor d(319) xor d(318) xor d(313) xor d(310) xor d(309) xor d(308) xor d(307) xor d(306) xor d(303) xor d(301) xor d(300) xor d(299) xor d(297) xor d(296) xor d(289) xor d(288) xor d(287) xor d(286) xor d(283) xor d(282) xor d(281) xor d(280) xor d(279) xor d(275) xor d(274) xor d(270) xor d(268) xor d(267) xor d(266) xor d(262) xor d(261) xor d(259) xor d(257) xor d(255) xor d(253) xor d(252) xor d(251) xor d(249) xor d(246) xor d(245) xor d(244) xor d(242) xor d(241) xor d(237) xor d(234) xor d(232) xor d(231) xor d(229) xor d(224) xor d(223) xor d(222) xor d(220) xor d(219) xor d(217) xor d(214) xor d(213) xor d(207) xor d(206) xor d(204) xor d(202) xor d(199) xor d(197) xor d(193) xor d(192) xor d(191) xor d(190) xor d(189) xor d(187) xor d(184) xor d(183) xor d(182) xor d(179) xor d(177) xor d(176) xor d(175) xor d(172) xor d(171) xor d(168) xor d(167) xor d(164) xor d(163) xor d(162) xor d(159) xor d(156) xor d(153) xor d(152) xor d(151) xor d(149) xor d(148) xor d(147) xor d(145) xor d(143) xor d(142) xor d(141) xor d(140) xor d(138) xor d(135) xor d(133) xor d(131) xor d(129) xor d(126) xor d(124) xor d(122) xor d(119) xor d(116) xor d(111) xor d(110) xor d(109) xor d(108) xor d(106) xor d(105) xor d(104) xor d(103) xor d(98) xor d(97) xor d(95) xor d(93) xor d(87) xor d(80) xor d(79) xor d(77) xor d(76) xor d(75) xor d(74) xor d(71) xor d(69) xor d(68) xor d(60) xor d(58) xor d(57) xor d(56) xor d(54) xor d(52) xor d(51) xor d(50) xor d(47) xor d(46) xor d(45) xor d(43) xor d(42) xor d(41) xor d(39) xor d(37) xor d(34) xor d(32) xor d(29) xor d(28) xor d(25) xor d(24) xor d(23) xor d(22) xor d(21) xor d(16) xor d(15) xor d(10) xor d(8) xor d(7) xor d(5) xor d(3) xor d(2) xor d(0) xor c(1) xor c(2) xor c(3) xor c(6) xor c(7) xor c(8) xor c(10) xor c(13) xor c(14) xor c(16) xor c(17) xor c(19) xor c(21) xor c(22) xor c(26) xor c(29) xor c(30) xor c(31);
    newcrc(8) := d(508) xor d(506) xor d(503) xor d(501) xor d(498) xor d(497) xor d(493) xor d(492) xor d(490) xor d(487) xor d(486) xor d(484) xor d(481) xor d(480) xor d(479) xor d(478) xor d(477) xor d(473) xor d(470) xor d(468) xor d(466) xor d(465) xor d(464) xor d(463) xor d(462) xor d(460) xor d(458) xor d(455) xor d(453) xor d(451) xor d(450) xor d(447) xor d(444) xor d(441) xor d(435) xor d(433) xor d(432) xor d(431) xor d(429) xor d(426) xor d(424) xor d(423) xor d(422) xor d(418) xor d(417) xor d(415) xor d(414) xor d(412) xor d(410) xor d(409) xor d(408) xor d(403) xor d(402) xor d(401) xor d(400) xor d(396) xor d(393) xor d(390) xor d(389) xor d(388) xor d(387) xor d(384) xor d(383) xor d(381) xor d(380) xor d(379) xor d(378) xor d(377) xor d(374) xor d(373) xor d(369) xor d(367) xor d(366) xor d(364) xor d(362) xor d(361) xor d(360) xor d(359) xor d(357) xor d(356) xor d(355) xor d(354) xor d(349) xor d(345) xor d(337) xor d(336) xor d(332) xor d(329) xor d(328) xor d(325) xor d(323) xor d(322) xor d(321) xor d(318) xor d(317) xor d(315) xor d(314) xor d(312) xor d(311) xor d(308) xor d(307) xor d(305) xor d(304) xor d(303) xor d(301) xor d(299) xor d(296) xor d(295) xor d(294) xor d(292) xor d(289) xor d(286) xor d(284) xor d(282) xor d(281) xor d(280) xor d(279) xor d(277) xor d(275) xor d(274) xor d(273) xor d(271) xor d(267) xor d(265) xor d(264) xor d(263) xor d(262) xor d(261) xor d(260) xor d(259) xor d(258) xor d(257) xor d(256) xor d(255) xor d(254) xor d(253) xor d(250) xor d(248) xor d(247) xor d(246) xor d(245) xor d(242) xor d(238) xor d(237) xor d(235) xor d(234) xor d(233) xor d(232) xor d(228) xor d(227) xor d(226) xor d(225) xor d(223) xor d(221) xor d(220) xor d(218) xor d(216) xor d(215) xor d(212) xor d(210) xor d(209) xor d(205) xor d(202) xor d(201) xor d(200) xor d(199) xor d(197) xor d(186) xor d(185) xor d(184) xor d(182) xor d(180) xor d(178) xor d(177) xor d(176) xor d(173) xor d(171) xor d(170) xor d(168) xor d(167) xor d(166) xor d(165) xor d(164) xor d(163) xor d(162) xor d(161) xor d(160) xor d(158) xor d(157) xor d(156) xor d(155) xor d(154) xor d(153) xor d(152) xor d(151) xor d(150) xor d(148) xor d(146) xor d(142) xor d(141) xor d(139) xor d(137) xor d(135) xor d(130) xor d(128) xor d(126) xor d(120) xor d(119) xor d(118) xor d(116) xor d(114) xor d(113) xor d(112) xor d(109) xor d(107) xor d(105) xor d(103) xor d(101) xor d(97) xor d(95) xor d(88) xor d(87) xor d(85) xor d(84) xor d(83) xor d(82) xor d(80) xor d(79) xor d(78) xor d(77) xor d(76) xor d(75) xor d(73) xor d(70) xor d(69) xor d(68) xor d(67) xor d(66) xor d(65) xor d(63) xor d(60) xor d(59) xor d(57) xor d(54) xor d(52) xor d(51) xor d(50) xor d(46) xor d(45) xor d(43) xor d(42) xor d(40) xor d(38) xor d(37) xor d(35) xor d(34) xor d(33) xor d(32) xor d(31) xor d(28) xor d(23) xor d(22) xor d(17) xor d(12) xor d(11) xor d(10) xor d(8) xor d(4) xor d(3) xor d(1) xor d(0) xor c(0) xor c(1) xor c(4) xor c(6) xor c(7) xor c(10) xor c(12) xor c(13) xor c(17) xor c(18) xor c(21) xor c(23) xor c(26) xor c(28);
    newcrc(9) := d(509) xor d(507) xor d(504) xor d(502) xor d(499) xor d(498) xor d(494) xor d(493) xor d(491) xor d(488) xor d(487) xor d(485) xor d(482) xor d(481) xor d(480) xor d(479) xor d(478) xor d(474) xor d(471) xor d(469) xor d(467) xor d(466) xor d(465) xor d(464) xor d(463) xor d(461) xor d(459) xor d(456) xor d(454) xor d(452) xor d(451) xor d(448) xor d(445) xor d(442) xor d(436) xor d(434) xor d(433) xor d(432) xor d(430) xor d(427) xor d(425) xor d(424) xor d(423) xor d(419) xor d(418) xor d(416) xor d(415) xor d(413) xor d(411) xor d(410) xor d(409) xor d(404) xor d(403) xor d(402) xor d(401) xor d(397) xor d(394) xor d(391) xor d(390) xor d(389) xor d(388) xor d(385) xor d(384) xor d(382) xor d(381) xor d(380) xor d(379) xor d(378) xor d(375) xor d(374) xor d(370) xor d(368) xor d(367) xor d(365) xor d(363) xor d(362) xor d(361) xor d(360) xor d(358) xor d(357) xor d(356) xor d(355) xor d(350) xor d(346) xor d(338) xor d(337) xor d(333) xor d(330) xor d(329) xor d(326) xor d(324) xor d(323) xor d(322) xor d(319) xor d(318) xor d(316) xor d(315) xor d(313) xor d(312) xor d(309) xor d(308) xor d(306) xor d(305) xor d(304) xor d(302) xor d(300) xor d(297) xor d(296) xor d(295) xor d(293) xor d(290) xor d(287) xor d(285) xor d(283) xor d(282) xor d(281) xor d(280) xor d(278) xor d(276) xor d(275) xor d(274) xor d(272) xor d(268) xor d(266) xor d(265) xor d(264) xor d(263) xor d(262) xor d(261) xor d(260) xor d(259) xor d(258) xor d(257) xor d(256) xor d(255) xor d(254) xor d(251) xor d(249) xor d(248) xor d(247) xor d(246) xor d(243) xor d(239) xor d(238) xor d(236) xor d(235) xor d(234) xor d(233) xor d(229) xor d(228) xor d(227) xor d(226) xor d(224) xor d(222) xor d(221) xor d(219) xor d(217) xor d(216) xor d(213) xor d(211) xor d(210) xor d(206) xor d(203) xor d(202) xor d(201) xor d(200) xor d(198) xor d(187) xor d(186) xor d(185) xor d(183) xor d(181) xor d(179) xor d(178) xor d(177) xor d(174) xor d(172) xor d(171) xor d(169) xor d(168) xor d(167) xor d(166) xor d(165) xor d(164) xor d(163) xor d(162) xor d(161) xor d(159) xor d(158) xor d(157) xor d(156) xor d(155) xor d(154) xor d(153) xor d(152) xor d(151) xor d(149) xor d(147) xor d(143) xor d(142) xor d(140) xor d(138) xor d(136) xor d(131) xor d(129) xor d(127) xor d(121) xor d(120) xor d(119) xor d(117) xor d(115) xor d(114) xor d(113) xor d(110) xor d(108) xor d(106) xor d(104) xor d(102) xor d(98) xor d(96) xor d(89) xor d(88) xor d(86) xor d(85) xor d(84) xor d(83) xor d(81) xor d(80) xor d(79) xor d(78) xor d(77) xor d(76) xor d(74) xor d(71) xor d(70) xor d(69) xor d(68) xor d(67) xor d(66) xor d(64) xor d(61) xor d(60) xor d(58) xor d(55) xor d(53) xor d(52) xor d(51) xor d(47) xor d(46) xor d(44) xor d(43) xor d(41) xor d(39) xor d(38) xor d(36) xor d(35) xor d(34) xor d(33) xor d(32) xor d(29) xor d(24) xor d(23) xor d(18) xor d(13) xor d(12) xor d(11) xor d(9) xor d(5) xor d(4) xor d(2) xor d(1) xor c(0) xor c(1) xor c(2) xor c(5) xor c(7) xor c(8) xor c(11) xor c(13) xor c(14) xor c(18) xor c(19) xor c(22) xor c(24) xor c(27) xor c(29);
    newcrc(10) := d(511) xor d(507) xor d(506) xor d(505) xor d(503) xor d(502) xor d(501) xor d(499) xor d(493) xor d(491) xor d(490) xor d(477) xor d(476) xor d(475) xor d(467) xor d(466) xor d(461) xor d(460) xor d(458) xor d(457) xor d(455) xor d(453) xor d(450) xor d(448) xor d(446) xor d(444) xor d(443) xor d(436) xor d(435) xor d(431) xor d(428) xor d(426) xor d(425) xor d(422) xor d(420) xor d(418) xor d(417) xor d(411) xor d(410) xor d(409) xor d(408) xor d(407) xor d(403) xor d(402) xor d(400) xor d(399) xor d(396) xor d(395) xor d(393) xor d(389) xor d(388) xor d(387) xor d(385) xor d(383) xor d(382) xor d(380) xor d(379) xor d(378) xor d(375) xor d(374) xor d(372) xor d(371) xor d(364) xor d(361) xor d(356) xor d(353) xor d(351) xor d(349) xor d(348) xor d(345) xor d(344) xor d(342) xor d(341) xor d(337) xor d(335) xor d(333) xor d(331) xor d(330) xor d(328) xor d(325) xor d(324) xor d(323) xor d(322) xor d(321) xor d(318) xor d(316) xor d(315) xor d(314) xor d(313) xor d(312) xor d(307) xor d(306) xor d(302) xor d(301) xor d(300) xor d(299) xor d(295) xor d(292) xor d(291) xor d(290) xor d(287) xor d(284) xor d(282) xor d(281) xor d(275) xor d(274) xor d(268) xor d(267) xor d(266) xor d(263) xor d(262) xor d(260) xor d(258) xor d(256) xor d(250) xor d(249) xor d(247) xor d(244) xor d(243) xor d(240) xor d(239) xor d(236) xor d(235) xor d(229) xor d(226) xor d(225) xor d(224) xor d(223) xor d(222) xor d(220) xor d(218) xor d(217) xor d(216) xor d(211) xor d(210) xor d(209) xor d(208) xor d(204) xor d(198) xor d(197) xor d(194) xor d(193) xor d(192) xor d(191) xor d(190) xor d(187) xor d(184) xor d(183) xor d(180) xor d(179) xor d(178) xor d(175) xor d(173) xor d(171) xor d(168) xor d(165) xor d(164) xor d(163) xor d(161) xor d(160) xor d(159) xor d(157) xor d(154) xor d(153) xor d(152) xor d(151) xor d(150) xor d(149) xor d(148) xor d(141) xor d(139) xor d(136) xor d(135) xor d(134) xor d(130) xor d(127) xor d(126) xor d(125) xor d(123) xor d(122) xor d(121) xor d(120) xor d(119) xor d(117) xor d(115) xor d(113) xor d(110) xor d(109) xor d(107) xor d(106) xor d(105) xor d(104) xor d(101) xor d(98) xor d(96) xor d(95) xor d(94) xor d(90) xor d(89) xor d(86) xor d(83) xor d(80) xor d(78) xor d(77) xor d(75) xor d(73) xor d(71) xor d(70) xor d(69) xor d(66) xor d(63) xor d(62) xor d(60) xor d(59) xor d(58) xor d(56) xor d(55) xor d(52) xor d(50) xor d(42) xor d(40) xor d(39) xor d(36) xor d(35) xor d(33) xor d(32) xor d(31) xor d(29) xor d(28) xor d(26) xor d(19) xor d(16) xor d(14) xor d(13) xor d(9) xor d(5) xor d(3) xor d(2) xor d(0) xor c(10) xor c(11) xor c(13) xor c(19) xor c(21) xor c(22) xor c(23) xor c(25) xor c(26) xor c(27) xor c(31);
    newcrc(11) := d(511) xor d(510) xor d(504) xor d(503) xor d(501) xor d(495) xor d(493) xor d(490) xor d(489) xor d(488) xor d(486) xor d(483) xor d(482) xor d(481) xor d(480) xor d(479) xor d(478) xor d(472) xor d(470) xor d(467) xor d(465) xor d(464) xor d(459) xor d(456) xor d(454) xor d(452) xor d(451) xor d(450) xor d(448) xor d(447) xor d(445) xor d(434) xor d(433) xor d(432) xor d(429) xor d(427) xor d(426) xor d(424) xor d(423) xor d(422) xor d(421) xor d(416) xor d(414) xor d(411) xor d(410) xor d(407) xor d(405) xor d(403) xor d(401) xor d(399) xor d(398) xor d(397) xor d(394) xor d(393) xor d(392) xor d(391) xor d(389) xor d(387) xor d(384) xor d(383) xor d(380) xor d(379) xor d(378) xor d(375) xor d(374) xor d(373) xor d(369) xor d(368) xor d(366) xor d(365) xor d(363) xor d(359) xor d(358) xor d(354) xor d(353) xor d(352) xor d(350) xor d(348) xor d(347) xor d(346) xor d(344) xor d(343) xor d(341) xor d(339) xor d(337) xor d(336) xor d(335) xor d(333) xor d(332) xor d(331) xor d(329) xor d(328) xor d(327) xor d(326) xor d(325) xor d(324) xor d(323) xor d(321) xor d(320) xor d(318) xor d(316) xor d(314) xor d(313) xor d(312) xor d(310) xor d(309) xor d(308) xor d(307) xor d(305) xor d(301) xor d(299) xor d(298) xor d(297) xor d(295) xor d(294) xor d(293) xor d(291) xor d(290) xor d(287) xor d(286) xor d(285) xor d(282) xor d(279) xor d(277) xor d(275) xor d(274) xor d(273) xor d(267) xor d(265) xor d(263) xor d(255) xor d(252) xor d(251) xor d(250) xor d(245) xor d(244) xor d(243) xor d(241) xor d(240) xor d(236) xor d(234) xor d(228) xor d(225) xor d(223) xor d(221) xor d(219) xor d(218) xor d(217) xor d(216) xor d(214) xor d(211) xor d(208) xor d(207) xor d(205) xor d(203) xor d(202) xor d(201) xor d(197) xor d(195) xor d(190) xor d(186) xor d(185) xor d(184) xor d(183) xor d(182) xor d(181) xor d(180) xor d(179) xor d(176) xor d(174) xor d(171) xor d(170) xor d(167) xor d(165) xor d(164) xor d(160) xor d(156) xor d(154) xor d(153) xor d(152) xor d(150) xor d(144) xor d(143) xor d(142) xor d(140) xor d(134) xor d(132) xor d(131) xor d(125) xor d(124) xor d(122) xor d(121) xor d(120) xor d(119) xor d(117) xor d(113) xor d(108) xor d(107) xor d(105) xor d(104) xor d(103) xor d(102) xor d(101) xor d(98) xor d(94) xor d(91) xor d(90) xor d(85) xor d(83) xor d(82) xor d(78) xor d(76) xor d(74) xor d(73) xor d(71) xor d(70) xor d(68) xor d(66) xor d(65) xor d(64) xor d(59) xor d(58) xor d(57) xor d(56) xor d(55) xor d(54) xor d(51) xor d(50) xor d(48) xor d(47) xor d(45) xor d(44) xor d(43) xor d(41) xor d(40) xor d(36) xor d(33) xor d(31) xor d(28) xor d(27) xor d(26) xor d(25) xor d(24) xor d(20) xor d(17) xor d(16) xor d(15) xor d(14) xor d(12) xor d(9) xor d(4) xor d(3) xor d(1) xor d(0) xor c(0) xor c(1) xor c(2) xor c(3) xor c(6) xor c(8) xor c(9) xor c(10) xor c(13) xor c(15) xor c(21) xor c(23) xor c(24) xor c(30) xor c(31);
    newcrc(12) := d(510) xor d(508) xor d(507) xor d(506) xor d(505) xor d(504) xor d(501) xor d(500) xor d(496) xor d(495) xor d(493) xor d(492) xor d(488) xor d(487) xor d(486) xor d(484) xor d(477) xor d(476) xor d(473) xor d(472) xor d(471) xor d(470) xor d(466) xor d(464) xor d(462) xor d(461) xor d(460) xor d(458) xor d(457) xor d(455) xor d(453) xor d(451) xor d(450) xor d(446) xor d(444) xor d(437) xor d(436) xor d(435) xor d(430) xor d(428) xor d(427) xor d(425) xor d(423) xor d(419) xor d(418) xor d(417) xor d(416) xor d(415) xor d(414) xor d(411) xor d(409) xor d(407) xor d(406) xor d(405) xor d(402) xor d(396) xor d(395) xor d(394) xor d(391) xor d(387) xor d(386) xor d(385) xor d(384) xor d(380) xor d(379) xor d(378) xor d(375) xor d(372) xor d(370) xor d(368) xor d(367) xor d(364) xor d(363) xor d(362) xor d(360) xor d(358) xor d(357) xor d(355) xor d(354) xor d(351) xor d(341) xor d(340) xor d(339) xor d(336) xor d(335) xor d(332) xor d(330) xor d(329) xor d(326) xor d(325) xor d(324) xor d(320) xor d(318) xor d(314) xor d(313) xor d(312) xor d(311) xor d(308) xor d(306) xor d(305) xor d(303) xor d(297) xor d(291) xor d(290) xor d(280) xor d(279) xor d(278) xor d(277) xor d(275) xor d(273) xor d(269) xor d(266) xor d(265) xor d(261) xor d(259) xor d(257) xor d(256) xor d(255) xor d(253) xor d(251) xor d(248) xor d(246) xor d(245) xor d(244) xor d(243) xor d(242) xor d(241) xor d(235) xor d(234) xor d(230) xor d(229) xor d(228) xor d(227) xor d(222) xor d(220) xor d(219) xor d(218) xor d(217) xor d(216) xor d(215) xor d(214) xor d(210) xor d(207) xor d(206) xor d(204) xor d(201) xor d(199) xor d(197) xor d(196) xor d(194) xor d(193) xor d(192) xor d(190) xor d(188) xor d(187) xor d(185) xor d(184) xor d(181) xor d(180) xor d(177) xor d(175) xor d(170) xor d(169) xor d(168) xor d(167) xor d(165) xor d(162) xor d(158) xor d(157) xor d(156) xor d(154) xor d(153) xor d(149) xor d(145) xor d(141) xor d(137) xor d(136) xor d(134) xor d(133) xor d(128) xor d(127) xor d(122) xor d(121) xor d(120) xor d(119) xor d(117) xor d(116) xor d(113) xor d(111) xor d(110) xor d(109) xor d(108) xor d(105) xor d(102) xor d(101) xor d(98) xor d(97) xor d(96) xor d(94) xor d(92) xor d(91) xor d(87) xor d(86) xor d(85) xor d(82) xor d(81) xor d(77) xor d(75) xor d(74) xor d(73) xor d(71) xor d(69) xor d(68) xor d(63) xor d(61) xor d(59) xor d(57) xor d(56) xor d(54) xor d(53) xor d(52) xor d(51) xor d(50) xor d(49) xor d(47) xor d(46) xor d(42) xor d(41) xor d(31) xor d(30) xor d(27) xor d(24) xor d(21) xor d(18) xor d(17) xor d(15) xor d(13) xor d(12) xor d(9) xor d(6) xor d(5) xor d(4) xor d(2) xor d(1) xor d(0) xor c(4) xor c(6) xor c(7) xor c(8) xor c(12) xor c(13) xor c(15) xor c(16) xor c(20) xor c(21) xor c(24) xor c(25) xor c(26) xor c(27) xor c(28) xor c(30);
    newcrc(13) := d(511) xor d(509) xor d(508) xor d(507) xor d(506) xor d(505) xor d(502) xor d(501) xor d(497) xor d(496) xor d(494) xor d(493) xor d(489) xor d(488) xor d(487) xor d(485) xor d(478) xor d(477) xor d(474) xor d(473) xor d(472) xor d(471) xor d(467) xor d(465) xor d(463) xor d(462) xor d(461) xor d(459) xor d(458) xor d(456) xor d(454) xor d(452) xor d(451) xor d(447) xor d(445) xor d(438) xor d(437) xor d(436) xor d(431) xor d(429) xor d(428) xor d(426) xor d(424) xor d(420) xor d(419) xor d(418) xor d(417) xor d(416) xor d(415) xor d(412) xor d(410) xor d(408) xor d(407) xor d(406) xor d(403) xor d(397) xor d(396) xor d(395) xor d(392) xor d(388) xor d(387) xor d(386) xor d(385) xor d(381) xor d(380) xor d(379) xor d(376) xor d(373) xor d(371) xor d(369) xor d(368) xor d(365) xor d(364) xor d(363) xor d(361) xor d(359) xor d(358) xor d(356) xor d(355) xor d(352) xor d(342) xor d(341) xor d(340) xor d(337) xor d(336) xor d(333) xor d(331) xor d(330) xor d(327) xor d(326) xor d(325) xor d(321) xor d(319) xor d(315) xor d(314) xor d(313) xor d(312) xor d(309) xor d(307) xor d(306) xor d(304) xor d(298) xor d(292) xor d(291) xor d(281) xor d(280) xor d(279) xor d(278) xor d(276) xor d(274) xor d(270) xor d(267) xor d(266) xor d(262) xor d(260) xor d(258) xor d(257) xor d(256) xor d(254) xor d(252) xor d(249) xor d(247) xor d(246) xor d(245) xor d(244) xor d(243) xor d(242) xor d(236) xor d(235) xor d(231) xor d(230) xor d(229) xor d(228) xor d(223) xor d(221) xor d(220) xor d(219) xor d(218) xor d(217) xor d(216) xor d(215) xor d(211) xor d(208) xor d(207) xor d(205) xor d(202) xor d(200) xor d(198) xor d(197) xor d(195) xor d(194) xor d(193) xor d(191) xor d(189) xor d(188) xor d(186) xor d(185) xor d(182) xor d(181) xor d(178) xor d(176) xor d(171) xor d(170) xor d(169) xor d(168) xor d(166) xor d(163) xor d(159) xor d(158) xor d(157) xor d(155) xor d(154) xor d(150) xor d(146) xor d(142) xor d(138) xor d(137) xor d(135) xor d(134) xor d(129) xor d(128) xor d(123) xor d(122) xor d(121) xor d(120) xor d(118) xor d(117) xor d(114) xor d(112) xor d(111) xor d(110) xor d(109) xor d(106) xor d(103) xor d(102) xor d(99) xor d(98) xor d(97) xor d(95) xor d(93) xor d(92) xor d(88) xor d(87) xor d(86) xor d(83) xor d(82) xor d(78) xor d(76) xor d(75) xor d(74) xor d(72) xor d(70) xor d(69) xor d(64) xor d(62) xor d(60) xor d(58) xor d(57) xor d(55) xor d(54) xor d(53) xor d(52) xor d(51) xor d(50) xor d(48) xor d(47) xor d(43) xor d(42) xor d(32) xor d(31) xor d(28) xor d(25) xor d(22) xor d(19) xor d(18) xor d(16) xor d(14) xor d(13) xor d(10) xor d(7) xor d(6) xor d(5) xor d(3) xor d(2) xor d(1) xor c(5) xor c(7) xor c(8) xor c(9) xor c(13) xor c(14) xor c(16) xor c(17) xor c(21) xor c(22) xor c(25) xor c(26) xor c(27) xor c(28) xor c(29) xor c(31);
    newcrc(14) := d(510) xor d(509) xor d(508) xor d(507) xor d(506) xor d(503) xor d(502) xor d(498) xor d(497) xor d(495) xor d(494) xor d(490) xor d(489) xor d(488) xor d(486) xor d(479) xor d(478) xor d(475) xor d(474) xor d(473) xor d(472) xor d(468) xor d(466) xor d(464) xor d(463) xor d(462) xor d(460) xor d(459) xor d(457) xor d(455) xor d(453) xor d(452) xor d(448) xor d(446) xor d(439) xor d(438) xor d(437) xor d(432) xor d(430) xor d(429) xor d(427) xor d(425) xor d(421) xor d(420) xor d(419) xor d(418) xor d(417) xor d(416) xor d(413) xor d(411) xor d(409) xor d(408) xor d(407) xor d(404) xor d(398) xor d(397) xor d(396) xor d(393) xor d(389) xor d(388) xor d(387) xor d(386) xor d(382) xor d(381) xor d(380) xor d(377) xor d(374) xor d(372) xor d(370) xor d(369) xor d(366) xor d(365) xor d(364) xor d(362) xor d(360) xor d(359) xor d(357) xor d(356) xor d(353) xor d(343) xor d(342) xor d(341) xor d(338) xor d(337) xor d(334) xor d(332) xor d(331) xor d(328) xor d(327) xor d(326) xor d(322) xor d(320) xor d(316) xor d(315) xor d(314) xor d(313) xor d(310) xor d(308) xor d(307) xor d(305) xor d(299) xor d(293) xor d(292) xor d(282) xor d(281) xor d(280) xor d(279) xor d(277) xor d(275) xor d(271) xor d(268) xor d(267) xor d(263) xor d(261) xor d(259) xor d(258) xor d(257) xor d(255) xor d(253) xor d(250) xor d(248) xor d(247) xor d(246) xor d(245) xor d(244) xor d(243) xor d(237) xor d(236) xor d(232) xor d(231) xor d(230) xor d(229) xor d(224) xor d(222) xor d(221) xor d(220) xor d(219) xor d(218) xor d(217) xor d(216) xor d(212) xor d(209) xor d(208) xor d(206) xor d(203) xor d(201) xor d(199) xor d(198) xor d(196) xor d(195) xor d(194) xor d(192) xor d(190) xor d(189) xor d(187) xor d(186) xor d(183) xor d(182) xor d(179) xor d(177) xor d(172) xor d(171) xor d(170) xor d(169) xor d(167) xor d(164) xor d(160) xor d(159) xor d(158) xor d(156) xor d(155) xor d(151) xor d(147) xor d(143) xor d(139) xor d(138) xor d(136) xor d(135) xor d(130) xor d(129) xor d(124) xor d(123) xor d(122) xor d(121) xor d(119) xor d(118) xor d(115) xor d(113) xor d(112) xor d(111) xor d(110) xor d(107) xor d(104) xor d(103) xor d(100) xor d(99) xor d(98) xor d(96) xor d(94) xor d(93) xor d(89) xor d(88) xor d(87) xor d(84) xor d(83) xor d(79) xor d(77) xor d(76) xor d(75) xor d(73) xor d(71) xor d(70) xor d(65) xor d(63) xor d(61) xor d(59) xor d(58) xor d(56) xor d(55) xor d(54) xor d(53) xor d(52) xor d(51) xor d(49) xor d(48) xor d(44) xor d(43) xor d(33) xor d(32) xor d(29) xor d(26) xor d(23) xor d(20) xor d(19) xor d(17) xor d(15) xor d(14) xor d(11) xor d(8) xor d(7) xor d(6) xor d(4) xor d(3) xor d(2) xor c(6) xor c(8) xor c(9) xor c(10) xor c(14) xor c(15) xor c(17) xor c(18) xor c(22) xor c(23) xor c(26) xor c(27) xor c(28) xor c(29) xor c(30);
    newcrc(15) := d(511) xor d(510) xor d(509) xor d(508) xor d(507) xor d(504) xor d(503) xor d(499) xor d(498) xor d(496) xor d(495) xor d(491) xor d(490) xor d(489) xor d(487) xor d(480) xor d(479) xor d(476) xor d(475) xor d(474) xor d(473) xor d(469) xor d(467) xor d(465) xor d(464) xor d(463) xor d(461) xor d(460) xor d(458) xor d(456) xor d(454) xor d(453) xor d(449) xor d(447) xor d(440) xor d(439) xor d(438) xor d(433) xor d(431) xor d(430) xor d(428) xor d(426) xor d(422) xor d(421) xor d(420) xor d(419) xor d(418) xor d(417) xor d(414) xor d(412) xor d(410) xor d(409) xor d(408) xor d(405) xor d(399) xor d(398) xor d(397) xor d(394) xor d(390) xor d(389) xor d(388) xor d(387) xor d(383) xor d(382) xor d(381) xor d(378) xor d(375) xor d(373) xor d(371) xor d(370) xor d(367) xor d(366) xor d(365) xor d(363) xor d(361) xor d(360) xor d(358) xor d(357) xor d(354) xor d(344) xor d(343) xor d(342) xor d(339) xor d(338) xor d(335) xor d(333) xor d(332) xor d(329) xor d(328) xor d(327) xor d(323) xor d(321) xor d(317) xor d(316) xor d(315) xor d(314) xor d(311) xor d(309) xor d(308) xor d(306) xor d(300) xor d(294) xor d(293) xor d(283) xor d(282) xor d(281) xor d(280) xor d(278) xor d(276) xor d(272) xor d(269) xor d(268) xor d(264) xor d(262) xor d(260) xor d(259) xor d(258) xor d(256) xor d(254) xor d(251) xor d(249) xor d(248) xor d(247) xor d(246) xor d(245) xor d(244) xor d(238) xor d(237) xor d(233) xor d(232) xor d(231) xor d(230) xor d(225) xor d(223) xor d(222) xor d(221) xor d(220) xor d(219) xor d(218) xor d(217) xor d(213) xor d(210) xor d(209) xor d(207) xor d(204) xor d(202) xor d(200) xor d(199) xor d(197) xor d(196) xor d(195) xor d(193) xor d(191) xor d(190) xor d(188) xor d(187) xor d(184) xor d(183) xor d(180) xor d(178) xor d(173) xor d(172) xor d(171) xor d(170) xor d(168) xor d(165) xor d(161) xor d(160) xor d(159) xor d(157) xor d(156) xor d(152) xor d(148) xor d(144) xor d(140) xor d(139) xor d(137) xor d(136) xor d(131) xor d(130) xor d(125) xor d(124) xor d(123) xor d(122) xor d(120) xor d(119) xor d(116) xor d(114) xor d(113) xor d(112) xor d(111) xor d(108) xor d(105) xor d(104) xor d(101) xor d(100) xor d(99) xor d(97) xor d(95) xor d(94) xor d(90) xor d(89) xor d(88) xor d(85) xor d(84) xor d(80) xor d(78) xor d(77) xor d(76) xor d(74) xor d(72) xor d(71) xor d(66) xor d(64) xor d(62) xor d(60) xor d(59) xor d(57) xor d(56) xor d(55) xor d(54) xor d(53) xor d(52) xor d(50) xor d(49) xor d(45) xor d(44) xor d(34) xor d(33) xor d(30) xor d(27) xor d(24) xor d(21) xor d(20) xor d(18) xor d(16) xor d(15) xor d(12) xor d(9) xor d(8) xor d(7) xor d(5) xor d(4) xor d(3) xor c(0) xor c(7) xor c(9) xor c(10) xor c(11) xor c(15) xor c(16) xor c(18) xor c(19) xor c(23) xor c(24) xor c(27) xor c(28) xor c(29) xor c(30) xor c(31);
    newcrc(16) := d(509) xor d(507) xor d(506) xor d(505) xor d(504) xor d(502) xor d(501) xor d(499) xor d(497) xor d(496) xor d(495) xor d(494) xor d(493) xor d(489) xor d(486) xor d(483) xor d(482) xor d(479) xor d(475) xor d(474) xor d(472) xor d(466) xor d(459) xor d(458) xor d(457) xor d(455) xor d(454) xor d(452) xor d(449) xor d(444) xor d(441) xor d(440) xor d(439) xor d(437) xor d(436) xor d(433) xor d(432) xor d(431) xor d(429) xor d(427) xor d(424) xor d(423) xor d(421) xor d(420) xor d(416) xor d(415) xor d(414) xor d(413) xor d(412) xor d(411) xor d(410) xor d(408) xor d(407) xor d(406) xor d(405) xor d(404) xor d(396) xor d(395) xor d(393) xor d(392) xor d(389) xor d(387) xor d(386) xor d(384) xor d(383) xor d(382) xor d(381) xor d(379) xor d(378) xor d(371) xor d(369) xor d(367) xor d(364) xor d(363) xor d(361) xor d(357) xor d(355) xor d(353) xor d(349) xor d(348) xor d(347) xor d(343) xor d(342) xor d(341) xor d(340) xor d(338) xor d(337) xor d(336) xor d(335) xor d(330) xor d(329) xor d(327) xor d(324) xor d(321) xor d(320) xor d(319) xor d(316) xor d(307) xor d(305) xor d(303) xor d(302) xor d(301) xor d(300) xor d(299) xor d(298) xor d(297) xor d(296) xor d(292) xor d(290) xor d(288) xor d(287) xor d(286) xor d(284) xor d(282) xor d(281) xor d(276) xor d(274) xor d(270) xor d(268) xor d(264) xor d(263) xor d(260) xor d(250) xor d(249) xor d(247) xor d(246) xor d(245) xor d(243) xor d(239) xor d(238) xor d(237) xor d(233) xor d(232) xor d(231) xor d(230) xor d(228) xor d(227) xor d(223) xor d(222) xor d(221) xor d(220) xor d(219) xor d(218) xor d(216) xor d(212) xor d(211) xor d(209) xor d(207) xor d(205) xor d(202) xor d(200) xor d(199) xor d(196) xor d(193) xor d(190) xor d(189) xor d(186) xor d(185) xor d(184) xor d(183) xor d(182) xor d(181) xor d(179) xor d(174) xor d(173) xor d(170) xor d(167) xor d(160) xor d(157) xor d(156) xor d(155) xor d(153) xor d(151) xor d(145) xor d(144) xor d(143) xor d(141) xor d(140) xor d(138) xor d(136) xor d(135) xor d(134) xor d(131) xor d(128) xor d(127) xor d(124) xor d(121) xor d(120) xor d(119) xor d(118) xor d(116) xor d(115) xor d(112) xor d(111) xor d(110) xor d(109) xor d(105) xor d(104) xor d(103) xor d(102) xor d(100) xor d(99) xor d(97) xor d(94) xor d(91) xor d(90) xor d(89) xor d(87) xor d(86) xor d(84) xor d(83) xor d(82) xor d(78) xor d(77) xor d(75) xor d(68) xor d(66) xor d(57) xor d(56) xor d(51) xor d(48) xor d(47) xor d(46) xor d(44) xor d(37) xor d(35) xor d(32) xor d(30) xor d(29) xor d(26) xor d(24) xor d(22) xor d(21) xor d(19) xor d(17) xor d(13) xor d(12) xor d(8) xor d(5) xor d(4) xor d(0) xor c(2) xor c(3) xor c(6) xor c(9) xor c(13) xor c(14) xor c(15) xor c(16) xor c(17) xor c(19) xor c(21) xor c(22) xor c(24) xor c(25) xor c(26) xor c(27) xor c(29);
    newcrc(17) := d(510) xor d(508) xor d(507) xor d(506) xor d(505) xor d(503) xor d(502) xor d(500) xor d(498) xor d(497) xor d(496) xor d(495) xor d(494) xor d(490) xor d(487) xor d(484) xor d(483) xor d(480) xor d(476) xor d(475) xor d(473) xor d(467) xor d(460) xor d(459) xor d(458) xor d(456) xor d(455) xor d(453) xor d(450) xor d(445) xor d(442) xor d(441) xor d(440) xor d(438) xor d(437) xor d(434) xor d(433) xor d(432) xor d(430) xor d(428) xor d(425) xor d(424) xor d(422) xor d(421) xor d(417) xor d(416) xor d(415) xor d(414) xor d(413) xor d(412) xor d(411) xor d(409) xor d(408) xor d(407) xor d(406) xor d(405) xor d(397) xor d(396) xor d(394) xor d(393) xor d(390) xor d(388) xor d(387) xor d(385) xor d(384) xor d(383) xor d(382) xor d(380) xor d(379) xor d(372) xor d(370) xor d(368) xor d(365) xor d(364) xor d(362) xor d(358) xor d(356) xor d(354) xor d(350) xor d(349) xor d(348) xor d(344) xor d(343) xor d(342) xor d(341) xor d(339) xor d(338) xor d(337) xor d(336) xor d(331) xor d(330) xor d(328) xor d(325) xor d(322) xor d(321) xor d(320) xor d(317) xor d(308) xor d(306) xor d(304) xor d(303) xor d(302) xor d(301) xor d(300) xor d(299) xor d(298) xor d(297) xor d(293) xor d(291) xor d(289) xor d(288) xor d(287) xor d(285) xor d(283) xor d(282) xor d(277) xor d(275) xor d(271) xor d(269) xor d(265) xor d(264) xor d(261) xor d(251) xor d(250) xor d(248) xor d(247) xor d(246) xor d(244) xor d(240) xor d(239) xor d(238) xor d(234) xor d(233) xor d(232) xor d(231) xor d(229) xor d(228) xor d(224) xor d(223) xor d(222) xor d(221) xor d(220) xor d(219) xor d(217) xor d(213) xor d(212) xor d(210) xor d(208) xor d(206) xor d(203) xor d(201) xor d(200) xor d(197) xor d(194) xor d(191) xor d(190) xor d(187) xor d(186) xor d(185) xor d(184) xor d(183) xor d(182) xor d(180) xor d(175) xor d(174) xor d(171) xor d(168) xor d(161) xor d(158) xor d(157) xor d(156) xor d(154) xor d(152) xor d(146) xor d(145) xor d(144) xor d(142) xor d(141) xor d(139) xor d(137) xor d(136) xor d(135) xor d(132) xor d(129) xor d(128) xor d(125) xor d(122) xor d(121) xor d(120) xor d(119) xor d(117) xor d(116) xor d(113) xor d(112) xor d(111) xor d(110) xor d(106) xor d(105) xor d(104) xor d(103) xor d(101) xor d(100) xor d(98) xor d(95) xor d(92) xor d(91) xor d(90) xor d(88) xor d(87) xor d(85) xor d(84) xor d(83) xor d(79) xor d(78) xor d(76) xor d(69) xor d(67) xor d(58) xor d(57) xor d(52) xor d(49) xor d(48) xor d(47) xor d(45) xor d(38) xor d(36) xor d(33) xor d(31) xor d(30) xor d(27) xor d(25) xor d(23) xor d(22) xor d(20) xor d(18) xor d(14) xor d(13) xor d(9) xor d(6) xor d(5) xor d(1) xor c(0) xor c(3) xor c(4) xor c(7) xor c(10) xor c(14) xor c(15) xor c(16) xor c(17) xor c(18) xor c(20) xor c(22) xor c(23) xor c(25) xor c(26) xor c(27) xor c(28) xor c(30);
    newcrc(18) := d(511) xor d(509) xor d(508) xor d(507) xor d(506) xor d(504) xor d(503) xor d(501) xor d(499) xor d(498) xor d(497) xor d(496) xor d(495) xor d(491) xor d(488) xor d(485) xor d(484) xor d(481) xor d(477) xor d(476) xor d(474) xor d(468) xor d(461) xor d(460) xor d(459) xor d(457) xor d(456) xor d(454) xor d(451) xor d(446) xor d(443) xor d(442) xor d(441) xor d(439) xor d(438) xor d(435) xor d(434) xor d(433) xor d(431) xor d(429) xor d(426) xor d(425) xor d(423) xor d(422) xor d(418) xor d(417) xor d(416) xor d(415) xor d(414) xor d(413) xor d(412) xor d(410) xor d(409) xor d(408) xor d(407) xor d(406) xor d(398) xor d(397) xor d(395) xor d(394) xor d(391) xor d(389) xor d(388) xor d(386) xor d(385) xor d(384) xor d(383) xor d(381) xor d(380) xor d(373) xor d(371) xor d(369) xor d(366) xor d(365) xor d(363) xor d(359) xor d(357) xor d(355) xor d(351) xor d(350) xor d(349) xor d(345) xor d(344) xor d(343) xor d(342) xor d(340) xor d(339) xor d(338) xor d(337) xor d(332) xor d(331) xor d(329) xor d(326) xor d(323) xor d(322) xor d(321) xor d(318) xor d(309) xor d(307) xor d(305) xor d(304) xor d(303) xor d(302) xor d(301) xor d(300) xor d(299) xor d(298) xor d(294) xor d(292) xor d(290) xor d(289) xor d(288) xor d(286) xor d(284) xor d(283) xor d(278) xor d(276) xor d(272) xor d(270) xor d(266) xor d(265) xor d(262) xor d(252) xor d(251) xor d(249) xor d(248) xor d(247) xor d(245) xor d(241) xor d(240) xor d(239) xor d(235) xor d(234) xor d(233) xor d(232) xor d(230) xor d(229) xor d(225) xor d(224) xor d(223) xor d(222) xor d(221) xor d(220) xor d(218) xor d(214) xor d(213) xor d(211) xor d(209) xor d(207) xor d(204) xor d(202) xor d(201) xor d(198) xor d(195) xor d(192) xor d(191) xor d(188) xor d(187) xor d(186) xor d(185) xor d(184) xor d(183) xor d(181) xor d(176) xor d(175) xor d(172) xor d(169) xor d(162) xor d(159) xor d(158) xor d(157) xor d(155) xor d(153) xor d(147) xor d(146) xor d(145) xor d(143) xor d(142) xor d(140) xor d(138) xor d(137) xor d(136) xor d(133) xor d(130) xor d(129) xor d(126) xor d(123) xor d(122) xor d(121) xor d(120) xor d(118) xor d(117) xor d(114) xor d(113) xor d(112) xor d(111) xor d(107) xor d(106) xor d(105) xor d(104) xor d(102) xor d(101) xor d(99) xor d(96) xor d(93) xor d(92) xor d(91) xor d(89) xor d(88) xor d(86) xor d(85) xor d(84) xor d(80) xor d(79) xor d(77) xor d(70) xor d(68) xor d(59) xor d(58) xor d(53) xor d(50) xor d(49) xor d(48) xor d(46) xor d(39) xor d(37) xor d(34) xor d(32) xor d(31) xor d(28) xor d(26) xor d(24) xor d(23) xor d(21) xor d(19) xor d(15) xor d(14) xor d(10) xor d(7) xor d(6) xor d(2) xor c(1) xor c(4) xor c(5) xor c(8) xor c(11) xor c(15) xor c(16) xor c(17) xor c(18) xor c(19) xor c(21) xor c(23) xor c(24) xor c(26) xor c(27) xor c(28) xor c(29) xor c(31);
    newcrc(19) := d(510) xor d(509) xor d(508) xor d(507) xor d(505) xor d(504) xor d(502) xor d(500) xor d(499) xor d(498) xor d(497) xor d(496) xor d(492) xor d(489) xor d(486) xor d(485) xor d(482) xor d(478) xor d(477) xor d(475) xor d(469) xor d(462) xor d(461) xor d(460) xor d(458) xor d(457) xor d(455) xor d(452) xor d(447) xor d(444) xor d(443) xor d(442) xor d(440) xor d(439) xor d(436) xor d(435) xor d(434) xor d(432) xor d(430) xor d(427) xor d(426) xor d(424) xor d(423) xor d(419) xor d(418) xor d(417) xor d(416) xor d(415) xor d(414) xor d(413) xor d(411) xor d(410) xor d(409) xor d(408) xor d(407) xor d(399) xor d(398) xor d(396) xor d(395) xor d(392) xor d(390) xor d(389) xor d(387) xor d(386) xor d(385) xor d(384) xor d(382) xor d(381) xor d(374) xor d(372) xor d(370) xor d(367) xor d(366) xor d(364) xor d(360) xor d(358) xor d(356) xor d(352) xor d(351) xor d(350) xor d(346) xor d(345) xor d(344) xor d(343) xor d(341) xor d(340) xor d(339) xor d(338) xor d(333) xor d(332) xor d(330) xor d(327) xor d(324) xor d(323) xor d(322) xor d(319) xor d(310) xor d(308) xor d(306) xor d(305) xor d(304) xor d(303) xor d(302) xor d(301) xor d(300) xor d(299) xor d(295) xor d(293) xor d(291) xor d(290) xor d(289) xor d(287) xor d(285) xor d(284) xor d(279) xor d(277) xor d(273) xor d(271) xor d(267) xor d(266) xor d(263) xor d(253) xor d(252) xor d(250) xor d(249) xor d(248) xor d(246) xor d(242) xor d(241) xor d(240) xor d(236) xor d(235) xor d(234) xor d(233) xor d(231) xor d(230) xor d(226) xor d(225) xor d(224) xor d(223) xor d(222) xor d(221) xor d(219) xor d(215) xor d(214) xor d(212) xor d(210) xor d(208) xor d(205) xor d(203) xor d(202) xor d(199) xor d(196) xor d(193) xor d(192) xor d(189) xor d(188) xor d(187) xor d(186) xor d(185) xor d(184) xor d(182) xor d(177) xor d(176) xor d(173) xor d(170) xor d(163) xor d(160) xor d(159) xor d(158) xor d(156) xor d(154) xor d(148) xor d(147) xor d(146) xor d(144) xor d(143) xor d(141) xor d(139) xor d(138) xor d(137) xor d(134) xor d(131) xor d(130) xor d(127) xor d(124) xor d(123) xor d(122) xor d(121) xor d(119) xor d(118) xor d(115) xor d(114) xor d(113) xor d(112) xor d(108) xor d(107) xor d(106) xor d(105) xor d(103) xor d(102) xor d(100) xor d(97) xor d(94) xor d(93) xor d(92) xor d(90) xor d(89) xor d(87) xor d(86) xor d(85) xor d(81) xor d(80) xor d(78) xor d(71) xor d(69) xor d(60) xor d(59) xor d(54) xor d(51) xor d(50) xor d(49) xor d(47) xor d(40) xor d(38) xor d(35) xor d(33) xor d(32) xor d(29) xor d(27) xor d(25) xor d(24) xor d(22) xor d(20) xor d(16) xor d(15) xor d(11) xor d(8) xor d(7) xor d(3) xor c(2) xor c(5) xor c(6) xor c(9) xor c(12) xor c(16) xor c(17) xor c(18) xor c(19) xor c(20) xor c(22) xor c(24) xor c(25) xor c(27) xor c(28) xor c(29) xor c(30);
    newcrc(20) := d(511) xor d(510) xor d(509) xor d(508) xor d(506) xor d(505) xor d(503) xor d(501) xor d(500) xor d(499) xor d(498) xor d(497) xor d(493) xor d(490) xor d(487) xor d(486) xor d(483) xor d(479) xor d(478) xor d(476) xor d(470) xor d(463) xor d(462) xor d(461) xor d(459) xor d(458) xor d(456) xor d(453) xor d(448) xor d(445) xor d(444) xor d(443) xor d(441) xor d(440) xor d(437) xor d(436) xor d(435) xor d(433) xor d(431) xor d(428) xor d(427) xor d(425) xor d(424) xor d(420) xor d(419) xor d(418) xor d(417) xor d(416) xor d(415) xor d(414) xor d(412) xor d(411) xor d(410) xor d(409) xor d(408) xor d(400) xor d(399) xor d(397) xor d(396) xor d(393) xor d(391) xor d(390) xor d(388) xor d(387) xor d(386) xor d(385) xor d(383) xor d(382) xor d(375) xor d(373) xor d(371) xor d(368) xor d(367) xor d(365) xor d(361) xor d(359) xor d(357) xor d(353) xor d(352) xor d(351) xor d(347) xor d(346) xor d(345) xor d(344) xor d(342) xor d(341) xor d(340) xor d(339) xor d(334) xor d(333) xor d(331) xor d(328) xor d(325) xor d(324) xor d(323) xor d(320) xor d(311) xor d(309) xor d(307) xor d(306) xor d(305) xor d(304) xor d(303) xor d(302) xor d(301) xor d(300) xor d(296) xor d(294) xor d(292) xor d(291) xor d(290) xor d(288) xor d(286) xor d(285) xor d(280) xor d(278) xor d(274) xor d(272) xor d(268) xor d(267) xor d(264) xor d(254) xor d(253) xor d(251) xor d(250) xor d(249) xor d(247) xor d(243) xor d(242) xor d(241) xor d(237) xor d(236) xor d(235) xor d(234) xor d(232) xor d(231) xor d(227) xor d(226) xor d(225) xor d(224) xor d(223) xor d(222) xor d(220) xor d(216) xor d(215) xor d(213) xor d(211) xor d(209) xor d(206) xor d(204) xor d(203) xor d(200) xor d(197) xor d(194) xor d(193) xor d(190) xor d(189) xor d(188) xor d(187) xor d(186) xor d(185) xor d(183) xor d(178) xor d(177) xor d(174) xor d(171) xor d(164) xor d(161) xor d(160) xor d(159) xor d(157) xor d(155) xor d(149) xor d(148) xor d(147) xor d(145) xor d(144) xor d(142) xor d(140) xor d(139) xor d(138) xor d(135) xor d(132) xor d(131) xor d(128) xor d(125) xor d(124) xor d(123) xor d(122) xor d(120) xor d(119) xor d(116) xor d(115) xor d(114) xor d(113) xor d(109) xor d(108) xor d(107) xor d(106) xor d(104) xor d(103) xor d(101) xor d(98) xor d(95) xor d(94) xor d(93) xor d(91) xor d(90) xor d(88) xor d(87) xor d(86) xor d(82) xor d(81) xor d(79) xor d(72) xor d(70) xor d(61) xor d(60) xor d(55) xor d(52) xor d(51) xor d(50) xor d(48) xor d(41) xor d(39) xor d(36) xor d(34) xor d(33) xor d(30) xor d(28) xor d(26) xor d(25) xor d(23) xor d(21) xor d(17) xor d(16) xor d(12) xor d(9) xor d(8) xor d(4) xor c(3) xor c(6) xor c(7) xor c(10) xor c(13) xor c(17) xor c(18) xor c(19) xor c(20) xor c(21) xor c(23) xor c(25) xor c(26) xor c(28) xor c(29) xor c(30) xor c(31);
    newcrc(21) := d(511) xor d(510) xor d(509) xor d(507) xor d(506) xor d(504) xor d(502) xor d(501) xor d(500) xor d(499) xor d(498) xor d(494) xor d(491) xor d(488) xor d(487) xor d(484) xor d(480) xor d(479) xor d(477) xor d(471) xor d(464) xor d(463) xor d(462) xor d(460) xor d(459) xor d(457) xor d(454) xor d(449) xor d(446) xor d(445) xor d(444) xor d(442) xor d(441) xor d(438) xor d(437) xor d(436) xor d(434) xor d(432) xor d(429) xor d(428) xor d(426) xor d(425) xor d(421) xor d(420) xor d(419) xor d(418) xor d(417) xor d(416) xor d(415) xor d(413) xor d(412) xor d(411) xor d(410) xor d(409) xor d(401) xor d(400) xor d(398) xor d(397) xor d(394) xor d(392) xor d(391) xor d(389) xor d(388) xor d(387) xor d(386) xor d(384) xor d(383) xor d(376) xor d(374) xor d(372) xor d(369) xor d(368) xor d(366) xor d(362) xor d(360) xor d(358) xor d(354) xor d(353) xor d(352) xor d(348) xor d(347) xor d(346) xor d(345) xor d(343) xor d(342) xor d(341) xor d(340) xor d(335) xor d(334) xor d(332) xor d(329) xor d(326) xor d(325) xor d(324) xor d(321) xor d(312) xor d(310) xor d(308) xor d(307) xor d(306) xor d(305) xor d(304) xor d(303) xor d(302) xor d(301) xor d(297) xor d(295) xor d(293) xor d(292) xor d(291) xor d(289) xor d(287) xor d(286) xor d(281) xor d(279) xor d(275) xor d(273) xor d(269) xor d(268) xor d(265) xor d(255) xor d(254) xor d(252) xor d(251) xor d(250) xor d(248) xor d(244) xor d(243) xor d(242) xor d(238) xor d(237) xor d(236) xor d(235) xor d(233) xor d(232) xor d(228) xor d(227) xor d(226) xor d(225) xor d(224) xor d(223) xor d(221) xor d(217) xor d(216) xor d(214) xor d(212) xor d(210) xor d(207) xor d(205) xor d(204) xor d(201) xor d(198) xor d(195) xor d(194) xor d(191) xor d(190) xor d(189) xor d(188) xor d(187) xor d(186) xor d(184) xor d(179) xor d(178) xor d(175) xor d(172) xor d(165) xor d(162) xor d(161) xor d(160) xor d(158) xor d(156) xor d(150) xor d(149) xor d(148) xor d(146) xor d(145) xor d(143) xor d(141) xor d(140) xor d(139) xor d(136) xor d(133) xor d(132) xor d(129) xor d(126) xor d(125) xor d(124) xor d(123) xor d(121) xor d(120) xor d(117) xor d(116) xor d(115) xor d(114) xor d(110) xor d(109) xor d(108) xor d(107) xor d(105) xor d(104) xor d(102) xor d(99) xor d(96) xor d(95) xor d(94) xor d(92) xor d(91) xor d(89) xor d(88) xor d(87) xor d(83) xor d(82) xor d(80) xor d(73) xor d(71) xor d(62) xor d(61) xor d(56) xor d(53) xor d(52) xor d(51) xor d(49) xor d(42) xor d(40) xor d(37) xor d(35) xor d(34) xor d(31) xor d(29) xor d(27) xor d(26) xor d(24) xor d(22) xor d(18) xor d(17) xor d(13) xor d(10) xor d(9) xor d(5) xor c(0) xor c(4) xor c(7) xor c(8) xor c(11) xor c(14) xor c(18) xor c(19) xor c(20) xor c(21) xor c(22) xor c(24) xor c(26) xor c(27) xor c(29) xor c(30) xor c(31);
    newcrc(22) := d(506) xor d(505) xor d(503) xor d(499) xor d(494) xor d(493) xor d(491) xor d(490) xor d(486) xor d(485) xor d(483) xor d(482) xor d(479) xor d(478) xor d(477) xor d(476) xor d(470) xor d(468) xor d(463) xor d(462) xor d(460) xor d(455) xor d(452) xor d(449) xor d(448) xor d(447) xor d(446) xor d(445) xor d(444) xor d(443) xor d(442) xor d(439) xor d(438) xor d(436) xor d(435) xor d(434) xor d(430) xor d(429) xor d(427) xor d(426) xor d(424) xor d(421) xor d(420) xor d(417) xor d(413) xor d(411) xor d(410) xor d(409) xor d(408) xor d(407) xor d(405) xor d(404) xor d(402) xor d(401) xor d(400) xor d(396) xor d(395) xor d(391) xor d(389) xor d(386) xor d(385) xor d(384) xor d(381) xor d(378) xor d(377) xor d(376) xor d(375) xor d(374) xor d(373) xor d(372) xor d(370) xor d(368) xor d(367) xor d(366) xor d(362) xor d(361) xor d(358) xor d(357) xor d(355) xor d(354) xor d(346) xor d(345) xor d(343) xor d(339) xor d(338) xor d(337) xor d(336) xor d(334) xor d(330) xor d(328) xor d(326) xor d(325) xor d(321) xor d(320) xor d(319) xor d(318) xor d(317) xor d(315) xor d(313) xor d(312) xor d(311) xor d(310) xor d(308) xor d(307) xor d(306) xor d(304) xor d(300) xor d(299) xor d(297) xor d(295) xor d(293) xor d(286) xor d(283) xor d(282) xor d(280) xor d(279) xor d(277) xor d(273) xor d(270) xor d(268) xor d(266) xor d(265) xor d(264) xor d(261) xor d(259) xor d(257) xor d(256) xor d(253) xor d(251) xor d(249) xor d(248) xor d(245) xor d(244) xor d(239) xor d(238) xor d(236) xor d(233) xor d(230) xor d(229) xor d(225) xor d(222) xor d(218) xor d(217) xor d(216) xor d(215) xor d(214) xor d(213) xor d(212) xor d(211) xor d(210) xor d(209) xor d(207) xor d(206) xor d(205) xor d(203) xor d(201) xor d(198) xor d(197) xor d(196) xor d(195) xor d(194) xor d(193) xor d(189) xor d(187) xor d(186) xor d(185) xor d(183) xor d(182) xor d(180) xor d(179) xor d(176) xor d(173) xor d(172) xor d(171) xor d(170) xor d(169) xor d(167) xor d(163) xor d(159) xor d(158) xor d(157) xor d(156) xor d(155) xor d(150) xor d(147) xor d(146) xor d(143) xor d(142) xor d(141) xor d(140) xor d(136) xor d(135) xor d(133) xor d(132) xor d(130) xor d(128) xor d(124) xor d(123) xor d(122) xor d(121) xor d(119) xor d(115) xor d(114) xor d(113) xor d(109) xor d(108) xor d(105) xor d(104) xor d(101) xor d(100) xor d(99) xor d(98) xor d(94) xor d(93) xor d(92) xor d(90) xor d(89) xor d(88) xor d(87) xor d(85) xor d(82) xor d(79) xor d(74) xor d(73) xor d(68) xor d(67) xor d(66) xor d(65) xor d(62) xor d(61) xor d(60) xor d(58) xor d(57) xor d(55) xor d(52) xor d(48) xor d(47) xor d(45) xor d(44) xor d(43) xor d(41) xor d(38) xor d(37) xor d(36) xor d(35) xor d(34) xor d(31) xor d(29) xor d(27) xor d(26) xor d(24) xor d(23) xor d(19) xor d(18) xor d(16) xor d(14) xor d(12) xor d(11) xor d(9) xor d(0) xor c(2) xor c(3) xor c(5) xor c(6) xor c(10) xor c(11) xor c(13) xor c(14) xor c(19) xor c(23) xor c(25) xor c(26);
    newcrc(23) := d(511) xor d(510) xor d(508) xor d(504) xor d(502) xor d(501) xor d(493) xor d(490) xor d(489) xor d(488) xor d(487) xor d(484) xor d(482) xor d(481) xor d(478) xor d(476) xor d(472) xor d(471) xor d(470) xor d(469) xor d(468) xor d(465) xor d(463) xor d(462) xor d(458) xor d(456) xor d(453) xor d(452) xor d(447) xor d(446) xor d(445) xor d(443) xor d(440) xor d(439) xor d(435) xor d(434) xor d(433) xor d(431) xor d(430) xor d(428) xor d(427) xor d(425) xor d(424) xor d(421) xor d(419) xor d(416) xor d(411) xor d(410) xor d(407) xor d(406) xor d(404) xor d(403) xor d(402) xor d(401) xor d(400) xor d(399) xor d(398) xor d(397) xor d(393) xor d(391) xor d(388) xor d(385) xor d(382) xor d(381) xor d(379) xor d(377) xor d(375) xor d(373) xor d(372) xor d(371) xor d(367) xor d(366) xor d(357) xor d(356) xor d(355) xor d(353) xor d(349) xor d(348) xor d(346) xor d(345) xor d(342) xor d(341) xor d(340) xor d(334) xor d(333) xor d(331) xor d(329) xor d(328) xor d(326) xor d(317) xor d(316) xor d(315) xor d(314) xor d(313) xor d(311) xor d(310) xor d(308) xor d(307) xor d(303) xor d(302) xor d(301) xor d(299) xor d(297) xor d(295) xor d(292) xor d(290) xor d(288) xor d(286) xor d(284) xor d(281) xor d(280) xor d(279) xor d(278) xor d(277) xor d(276) xor d(273) xor d(271) xor d(268) xor d(267) xor d(266) xor d(264) xor d(262) xor d(261) xor d(260) xor d(259) xor d(258) xor d(255) xor d(254) xor d(250) xor d(249) xor d(248) xor d(246) xor d(245) xor d(243) xor d(240) xor d(239) xor d(231) xor d(228) xor d(227) xor d(224) xor d(223) xor d(219) xor d(218) xor d(217) xor d(215) xor d(213) xor d(211) xor d(209) xor d(206) xor d(204) xor d(203) xor d(201) xor d(196) xor d(195) xor d(193) xor d(192) xor d(191) xor d(187) xor d(184) xor d(182) xor d(181) xor d(180) xor d(177) xor d(174) xor d(173) xor d(169) xor d(168) xor d(167) xor d(166) xor d(164) xor d(162) xor d(161) xor d(160) xor d(159) xor d(157) xor d(155) xor d(149) xor d(148) xor d(147) xor d(142) xor d(141) xor d(135) xor d(133) xor d(132) xor d(131) xor d(129) xor d(128) xor d(127) xor d(126) xor d(124) xor d(122) xor d(120) xor d(119) xor d(118) xor d(117) xor d(115) xor d(113) xor d(111) xor d(109) xor d(105) xor d(104) xor d(103) xor d(102) xor d(100) xor d(98) xor d(97) xor d(96) xor d(93) xor d(91) xor d(90) xor d(89) xor d(88) xor d(87) xor d(86) xor d(85) xor d(84) xor d(82) xor d(81) xor d(80) xor d(79) xor d(75) xor d(74) xor d(73) xor d(72) xor d(69) xor d(65) xor d(62) xor d(60) xor d(59) xor d(56) xor d(55) xor d(54) xor d(50) xor d(49) xor d(47) xor d(46) xor d(42) xor d(39) xor d(38) xor d(36) xor d(35) xor d(34) xor d(31) xor d(29) xor d(27) xor d(26) xor d(20) xor d(19) xor d(17) xor d(16) xor d(15) xor d(13) xor d(9) xor d(6) xor d(1) xor d(0) xor c(1) xor c(2) xor c(4) xor c(7) xor c(8) xor c(9) xor c(10) xor c(13) xor c(21) xor c(22) xor c(24) xor c(28) xor c(30) xor c(31);
    newcrc(24) := d(511) xor d(509) xor d(505) xor d(503) xor d(502) xor d(494) xor d(491) xor d(490) xor d(489) xor d(488) xor d(485) xor d(483) xor d(482) xor d(479) xor d(477) xor d(473) xor d(472) xor d(471) xor d(470) xor d(469) xor d(466) xor d(464) xor d(463) xor d(459) xor d(457) xor d(454) xor d(453) xor d(448) xor d(447) xor d(446) xor d(444) xor d(441) xor d(440) xor d(436) xor d(435) xor d(434) xor d(432) xor d(431) xor d(429) xor d(428) xor d(426) xor d(425) xor d(422) xor d(420) xor d(417) xor d(412) xor d(411) xor d(408) xor d(407) xor d(405) xor d(404) xor d(403) xor d(402) xor d(401) xor d(400) xor d(399) xor d(398) xor d(394) xor d(392) xor d(389) xor d(386) xor d(383) xor d(382) xor d(380) xor d(378) xor d(376) xor d(374) xor d(373) xor d(372) xor d(368) xor d(367) xor d(358) xor d(357) xor d(356) xor d(354) xor d(350) xor d(349) xor d(347) xor d(346) xor d(343) xor d(342) xor d(341) xor d(335) xor d(334) xor d(332) xor d(330) xor d(329) xor d(327) xor d(318) xor d(317) xor d(316) xor d(315) xor d(314) xor d(312) xor d(311) xor d(309) xor d(308) xor d(304) xor d(303) xor d(302) xor d(300) xor d(298) xor d(296) xor d(293) xor d(291) xor d(289) xor d(287) xor d(285) xor d(282) xor d(281) xor d(280) xor d(279) xor d(278) xor d(277) xor d(274) xor d(272) xor d(269) xor d(268) xor d(267) xor d(265) xor d(263) xor d(262) xor d(261) xor d(260) xor d(259) xor d(256) xor d(255) xor d(251) xor d(250) xor d(249) xor d(247) xor d(246) xor d(244) xor d(241) xor d(240) xor d(232) xor d(229) xor d(228) xor d(225) xor d(224) xor d(220) xor d(219) xor d(218) xor d(216) xor d(214) xor d(212) xor d(210) xor d(207) xor d(205) xor d(204) xor d(202) xor d(197) xor d(196) xor d(194) xor d(193) xor d(192) xor d(188) xor d(185) xor d(183) xor d(182) xor d(181) xor d(178) xor d(175) xor d(174) xor d(170) xor d(169) xor d(168) xor d(167) xor d(165) xor d(163) xor d(162) xor d(161) xor d(160) xor d(158) xor d(156) xor d(150) xor d(149) xor d(148) xor d(143) xor d(142) xor d(136) xor d(134) xor d(133) xor d(132) xor d(130) xor d(129) xor d(128) xor d(127) xor d(125) xor d(123) xor d(121) xor d(120) xor d(119) xor d(118) xor d(116) xor d(114) xor d(112) xor d(110) xor d(106) xor d(105) xor d(104) xor d(103) xor d(101) xor d(99) xor d(98) xor d(97) xor d(94) xor d(92) xor d(91) xor d(90) xor d(89) xor d(88) xor d(87) xor d(86) xor d(85) xor d(83) xor d(82) xor d(81) xor d(80) xor d(76) xor d(75) xor d(74) xor d(73) xor d(70) xor d(66) xor d(63) xor d(61) xor d(60) xor d(57) xor d(56) xor d(55) xor d(51) xor d(50) xor d(48) xor d(47) xor d(43) xor d(40) xor d(39) xor d(37) xor d(36) xor d(35) xor d(32) xor d(30) xor d(28) xor d(27) xor d(21) xor d(20) xor d(18) xor d(17) xor d(16) xor d(14) xor d(10) xor d(7) xor d(2) xor d(1) xor c(2) xor c(3) xor c(5) xor c(8) xor c(9) xor c(10) xor c(11) xor c(14) xor c(22) xor c(23) xor c(25) xor c(29) xor c(31);
    newcrc(25) := d(510) xor d(506) xor d(504) xor d(503) xor d(495) xor d(492) xor d(491) xor d(490) xor d(489) xor d(486) xor d(484) xor d(483) xor d(480) xor d(478) xor d(474) xor d(473) xor d(472) xor d(471) xor d(470) xor d(467) xor d(465) xor d(464) xor d(460) xor d(458) xor d(455) xor d(454) xor d(449) xor d(448) xor d(447) xor d(445) xor d(442) xor d(441) xor d(437) xor d(436) xor d(435) xor d(433) xor d(432) xor d(430) xor d(429) xor d(427) xor d(426) xor d(423) xor d(421) xor d(418) xor d(413) xor d(412) xor d(409) xor d(408) xor d(406) xor d(405) xor d(404) xor d(403) xor d(402) xor d(401) xor d(400) xor d(399) xor d(395) xor d(393) xor d(390) xor d(387) xor d(384) xor d(383) xor d(381) xor d(379) xor d(377) xor d(375) xor d(374) xor d(373) xor d(369) xor d(368) xor d(359) xor d(358) xor d(357) xor d(355) xor d(351) xor d(350) xor d(348) xor d(347) xor d(344) xor d(343) xor d(342) xor d(336) xor d(335) xor d(333) xor d(331) xor d(330) xor d(328) xor d(319) xor d(318) xor d(317) xor d(316) xor d(315) xor d(313) xor d(312) xor d(310) xor d(309) xor d(305) xor d(304) xor d(303) xor d(301) xor d(299) xor d(297) xor d(294) xor d(292) xor d(290) xor d(288) xor d(286) xor d(283) xor d(282) xor d(281) xor d(280) xor d(279) xor d(278) xor d(275) xor d(273) xor d(270) xor d(269) xor d(268) xor d(266) xor d(264) xor d(263) xor d(262) xor d(261) xor d(260) xor d(257) xor d(256) xor d(252) xor d(251) xor d(250) xor d(248) xor d(247) xor d(245) xor d(242) xor d(241) xor d(233) xor d(230) xor d(229) xor d(226) xor d(225) xor d(221) xor d(220) xor d(219) xor d(217) xor d(215) xor d(213) xor d(211) xor d(208) xor d(206) xor d(205) xor d(203) xor d(198) xor d(197) xor d(195) xor d(194) xor d(193) xor d(189) xor d(186) xor d(184) xor d(183) xor d(182) xor d(179) xor d(176) xor d(175) xor d(171) xor d(170) xor d(169) xor d(168) xor d(166) xor d(164) xor d(163) xor d(162) xor d(161) xor d(159) xor d(157) xor d(151) xor d(150) xor d(149) xor d(144) xor d(143) xor d(137) xor d(135) xor d(134) xor d(133) xor d(131) xor d(130) xor d(129) xor d(128) xor d(126) xor d(124) xor d(122) xor d(121) xor d(120) xor d(119) xor d(117) xor d(115) xor d(113) xor d(111) xor d(107) xor d(106) xor d(105) xor d(104) xor d(102) xor d(100) xor d(99) xor d(98) xor d(95) xor d(93) xor d(92) xor d(91) xor d(90) xor d(89) xor d(88) xor d(87) xor d(86) xor d(84) xor d(83) xor d(82) xor d(81) xor d(77) xor d(76) xor d(75) xor d(74) xor d(71) xor d(67) xor d(64) xor d(62) xor d(61) xor d(58) xor d(57) xor d(56) xor d(52) xor d(51) xor d(49) xor d(48) xor d(44) xor d(41) xor d(40) xor d(38) xor d(37) xor d(36) xor d(33) xor d(31) xor d(29) xor d(28) xor d(22) xor d(21) xor d(19) xor d(18) xor d(17) xor d(15) xor d(11) xor d(8) xor d(3) xor d(2) xor c(0) xor c(3) xor c(4) xor c(6) xor c(9) xor c(10) xor c(11) xor c(12) xor c(15) xor c(23) xor c(24) xor c(26) xor c(30);
    newcrc(26) := d(510) xor d(508) xor d(506) xor d(505) xor d(504) xor d(502) xor d(501) xor d(500) xor d(496) xor d(495) xor d(494) xor d(489) xor d(488) xor d(487) xor d(486) xor d(485) xor d(484) xor d(483) xor d(482) xor d(480) xor d(477) xor d(476) xor d(475) xor d(474) xor d(473) xor d(471) xor d(470) xor d(466) xor d(464) xor d(462) xor d(459) xor d(458) xor d(456) xor d(455) xor d(452) xor d(446) xor d(444) xor d(443) xor d(442) xor d(438) xor d(431) xor d(430) xor d(428) xor d(427) xor d(418) xor d(416) xor d(413) xor d(412) xor d(410) xor d(408) xor d(406) xor d(403) xor d(402) xor d(401) xor d(399) xor d(398) xor d(394) xor d(393) xor d(392) xor d(390) xor d(387) xor d(386) xor d(385) xor d(384) xor d(382) xor d(381) xor d(380) xor d(375) xor d(372) xor d(370) xor d(368) xor d(366) xor d(363) xor d(362) xor d(360) xor d(357) xor d(356) xor d(353) xor d(352) xor d(351) xor d(347) xor d(343) xor d(342) xor d(341) xor d(339) xor d(338) xor d(336) xor d(335) xor d(333) xor d(332) xor d(331) xor d(329) xor d(328) xor d(327) xor d(322) xor d(321) xor d(316) xor d(315) xor d(314) xor d(313) xor d(312) xor d(311) xor d(309) xor d(306) xor d(304) xor d(303) xor d(299) xor d(297) xor d(296) xor d(294) xor d(293) xor d(292) xor d(291) xor d(290) xor d(289) xor d(288) xor d(286) xor d(284) xor d(282) xor d(281) xor d(280) xor d(277) xor d(273) xor d(271) xor d(270) xor d(268) xor d(267) xor d(263) xor d(262) xor d(259) xor d(258) xor d(255) xor d(253) xor d(251) xor d(249) xor d(246) xor d(242) xor d(237) xor d(231) xor d(228) xor d(224) xor d(222) xor d(221) xor d(220) xor d(218) xor d(210) xor d(208) xor d(206) xor d(204) xor d(203) xor d(202) xor d(201) xor d(197) xor d(196) xor d(195) xor d(193) xor d(192) xor d(191) xor d(188) xor d(187) xor d(186) xor d(185) xor d(184) xor d(182) xor d(180) xor d(177) xor d(176) xor d(166) xor d(165) xor d(164) xor d(163) xor d(161) xor d(160) xor d(156) xor d(155) xor d(152) xor d(150) xor d(149) xor d(145) xor d(143) xor d(138) xor d(137) xor d(131) xor d(130) xor d(129) xor d(128) xor d(126) xor d(122) xor d(121) xor d(120) xor d(119) xor d(117) xor d(113) xor d(112) xor d(111) xor d(110) xor d(108) xor d(107) xor d(105) xor d(104) xor d(100) xor d(98) xor d(97) xor d(95) xor d(93) xor d(92) xor d(91) xor d(90) xor d(89) xor d(88) xor d(81) xor d(79) xor d(78) xor d(77) xor d(76) xor d(75) xor d(73) xor d(67) xor d(66) xor d(62) xor d(61) xor d(60) xor d(59) xor d(57) xor d(55) xor d(54) xor d(52) xor d(49) xor d(48) xor d(47) xor d(44) xor d(42) xor d(41) xor d(39) xor d(38) xor d(31) xor d(28) xor d(26) xor d(25) xor d(24) xor d(23) xor d(22) xor d(20) xor d(19) xor d(18) xor d(10) xor d(6) xor d(4) xor d(3) xor d(0) xor c(0) xor c(2) xor c(3) xor c(4) xor c(5) xor c(6) xor c(7) xor c(8) xor c(9) xor c(14) xor c(15) xor c(16) xor c(20) xor c(21) xor c(22) xor c(24) xor c(25) xor c(26) xor c(28) xor c(30);
    newcrc(27) := d(511) xor d(509) xor d(507) xor d(506) xor d(505) xor d(503) xor d(502) xor d(501) xor d(497) xor d(496) xor d(495) xor d(490) xor d(489) xor d(488) xor d(487) xor d(486) xor d(485) xor d(484) xor d(483) xor d(481) xor d(478) xor d(477) xor d(476) xor d(475) xor d(474) xor d(472) xor d(471) xor d(467) xor d(465) xor d(463) xor d(460) xor d(459) xor d(457) xor d(456) xor d(453) xor d(447) xor d(445) xor d(444) xor d(443) xor d(439) xor d(432) xor d(431) xor d(429) xor d(428) xor d(419) xor d(417) xor d(414) xor d(413) xor d(411) xor d(409) xor d(407) xor d(404) xor d(403) xor d(402) xor d(400) xor d(399) xor d(395) xor d(394) xor d(393) xor d(391) xor d(388) xor d(387) xor d(386) xor d(385) xor d(383) xor d(382) xor d(381) xor d(376) xor d(373) xor d(371) xor d(369) xor d(367) xor d(364) xor d(363) xor d(361) xor d(358) xor d(357) xor d(354) xor d(353) xor d(352) xor d(348) xor d(344) xor d(343) xor d(342) xor d(340) xor d(339) xor d(337) xor d(336) xor d(334) xor d(333) xor d(332) xor d(330) xor d(329) xor d(328) xor d(323) xor d(322) xor d(317) xor d(316) xor d(315) xor d(314) xor d(313) xor d(312) xor d(310) xor d(307) xor d(305) xor d(304) xor d(300) xor d(298) xor d(297) xor d(295) xor d(294) xor d(293) xor d(292) xor d(291) xor d(290) xor d(289) xor d(287) xor d(285) xor d(283) xor d(282) xor d(281) xor d(278) xor d(274) xor d(272) xor d(271) xor d(269) xor d(268) xor d(264) xor d(263) xor d(260) xor d(259) xor d(256) xor d(254) xor d(252) xor d(250) xor d(247) xor d(243) xor d(238) xor d(232) xor d(229) xor d(225) xor d(223) xor d(222) xor d(221) xor d(219) xor d(211) xor d(209) xor d(207) xor d(205) xor d(204) xor d(203) xor d(202) xor d(198) xor d(197) xor d(196) xor d(194) xor d(193) xor d(192) xor d(189) xor d(188) xor d(187) xor d(186) xor d(185) xor d(183) xor d(181) xor d(178) xor d(177) xor d(167) xor d(166) xor d(165) xor d(164) xor d(162) xor d(161) xor d(157) xor d(156) xor d(153) xor d(151) xor d(150) xor d(146) xor d(144) xor d(139) xor d(138) xor d(132) xor d(131) xor d(130) xor d(129) xor d(127) xor d(123) xor d(122) xor d(121) xor d(120) xor d(118) xor d(114) xor d(113) xor d(112) xor d(111) xor d(109) xor d(108) xor d(106) xor d(105) xor d(101) xor d(99) xor d(98) xor d(96) xor d(94) xor d(93) xor d(92) xor d(91) xor d(90) xor d(89) xor d(82) xor d(80) xor d(79) xor d(78) xor d(77) xor d(76) xor d(74) xor d(68) xor d(67) xor d(63) xor d(62) xor d(61) xor d(60) xor d(58) xor d(56) xor d(55) xor d(53) xor d(50) xor d(49) xor d(48) xor d(45) xor d(43) xor d(42) xor d(40) xor d(39) xor d(32) xor d(29) xor d(27) xor d(26) xor d(25) xor d(24) xor d(23) xor d(21) xor d(20) xor d(19) xor d(11) xor d(7) xor d(5) xor d(4) xor d(1) xor c(1) xor c(3) xor c(4) xor c(5) xor c(6) xor c(7) xor c(8) xor c(9) xor c(10) xor c(15) xor c(16) xor c(17) xor c(21) xor c(22) xor c(23) xor c(25) xor c(26) xor c(27) xor c(29) xor c(31);
    newcrc(28) := d(510) xor d(508) xor d(507) xor d(506) xor d(504) xor d(503) xor d(502) xor d(498) xor d(497) xor d(496) xor d(491) xor d(490) xor d(489) xor d(488) xor d(487) xor d(486) xor d(485) xor d(484) xor d(482) xor d(479) xor d(478) xor d(477) xor d(476) xor d(475) xor d(473) xor d(472) xor d(468) xor d(466) xor d(464) xor d(461) xor d(460) xor d(458) xor d(457) xor d(454) xor d(448) xor d(446) xor d(445) xor d(444) xor d(440) xor d(433) xor d(432) xor d(430) xor d(429) xor d(420) xor d(418) xor d(415) xor d(414) xor d(412) xor d(410) xor d(408) xor d(405) xor d(404) xor d(403) xor d(401) xor d(400) xor d(396) xor d(395) xor d(394) xor d(392) xor d(389) xor d(388) xor d(387) xor d(386) xor d(384) xor d(383) xor d(382) xor d(377) xor d(374) xor d(372) xor d(370) xor d(368) xor d(365) xor d(364) xor d(362) xor d(359) xor d(358) xor d(355) xor d(354) xor d(353) xor d(349) xor d(345) xor d(344) xor d(343) xor d(341) xor d(340) xor d(338) xor d(337) xor d(335) xor d(334) xor d(333) xor d(331) xor d(330) xor d(329) xor d(324) xor d(323) xor d(318) xor d(317) xor d(316) xor d(315) xor d(314) xor d(313) xor d(311) xor d(308) xor d(306) xor d(305) xor d(301) xor d(299) xor d(298) xor d(296) xor d(295) xor d(294) xor d(293) xor d(292) xor d(291) xor d(290) xor d(288) xor d(286) xor d(284) xor d(283) xor d(282) xor d(279) xor d(275) xor d(273) xor d(272) xor d(270) xor d(269) xor d(265) xor d(264) xor d(261) xor d(260) xor d(257) xor d(255) xor d(253) xor d(251) xor d(248) xor d(244) xor d(239) xor d(233) xor d(230) xor d(226) xor d(224) xor d(223) xor d(222) xor d(220) xor d(212) xor d(210) xor d(208) xor d(206) xor d(205) xor d(204) xor d(203) xor d(199) xor d(198) xor d(197) xor d(195) xor d(194) xor d(193) xor d(190) xor d(189) xor d(188) xor d(187) xor d(186) xor d(184) xor d(182) xor d(179) xor d(178) xor d(168) xor d(167) xor d(166) xor d(165) xor d(163) xor d(162) xor d(158) xor d(157) xor d(154) xor d(152) xor d(151) xor d(147) xor d(145) xor d(140) xor d(139) xor d(133) xor d(132) xor d(131) xor d(130) xor d(128) xor d(124) xor d(123) xor d(122) xor d(121) xor d(119) xor d(115) xor d(114) xor d(113) xor d(112) xor d(110) xor d(109) xor d(107) xor d(106) xor d(102) xor d(100) xor d(99) xor d(97) xor d(95) xor d(94) xor d(93) xor d(92) xor d(91) xor d(90) xor d(83) xor d(81) xor d(80) xor d(79) xor d(78) xor d(77) xor d(75) xor d(69) xor d(68) xor d(64) xor d(63) xor d(62) xor d(61) xor d(59) xor d(57) xor d(56) xor d(54) xor d(51) xor d(50) xor d(49) xor d(46) xor d(44) xor d(43) xor d(41) xor d(40) xor d(33) xor d(30) xor d(28) xor d(27) xor d(26) xor d(25) xor d(24) xor d(22) xor d(21) xor d(20) xor d(12) xor d(8) xor d(6) xor d(5) xor d(2) xor c(2) xor c(4) xor c(5) xor c(6) xor c(7) xor c(8) xor c(9) xor c(10) xor c(11) xor c(16) xor c(17) xor c(18) xor c(22) xor c(23) xor c(24) xor c(26) xor c(27) xor c(28) xor c(30);
    newcrc(29) := d(511) xor d(509) xor d(508) xor d(507) xor d(505) xor d(504) xor d(503) xor d(499) xor d(498) xor d(497) xor d(492) xor d(491) xor d(490) xor d(489) xor d(488) xor d(487) xor d(486) xor d(485) xor d(483) xor d(480) xor d(479) xor d(478) xor d(477) xor d(476) xor d(474) xor d(473) xor d(469) xor d(467) xor d(465) xor d(462) xor d(461) xor d(459) xor d(458) xor d(455) xor d(449) xor d(447) xor d(446) xor d(445) xor d(441) xor d(434) xor d(433) xor d(431) xor d(430) xor d(421) xor d(419) xor d(416) xor d(415) xor d(413) xor d(411) xor d(409) xor d(406) xor d(405) xor d(404) xor d(402) xor d(401) xor d(397) xor d(396) xor d(395) xor d(393) xor d(390) xor d(389) xor d(388) xor d(387) xor d(385) xor d(384) xor d(383) xor d(378) xor d(375) xor d(373) xor d(371) xor d(369) xor d(366) xor d(365) xor d(363) xor d(360) xor d(359) xor d(356) xor d(355) xor d(354) xor d(350) xor d(346) xor d(345) xor d(344) xor d(342) xor d(341) xor d(339) xor d(338) xor d(336) xor d(335) xor d(334) xor d(332) xor d(331) xor d(330) xor d(325) xor d(324) xor d(319) xor d(318) xor d(317) xor d(316) xor d(315) xor d(314) xor d(312) xor d(309) xor d(307) xor d(306) xor d(302) xor d(300) xor d(299) xor d(297) xor d(296) xor d(295) xor d(294) xor d(293) xor d(292) xor d(291) xor d(289) xor d(287) xor d(285) xor d(284) xor d(283) xor d(280) xor d(276) xor d(274) xor d(273) xor d(271) xor d(270) xor d(266) xor d(265) xor d(262) xor d(261) xor d(258) xor d(256) xor d(254) xor d(252) xor d(249) xor d(245) xor d(240) xor d(234) xor d(231) xor d(227) xor d(225) xor d(224) xor d(223) xor d(221) xor d(213) xor d(211) xor d(209) xor d(207) xor d(206) xor d(205) xor d(204) xor d(200) xor d(199) xor d(198) xor d(196) xor d(195) xor d(194) xor d(191) xor d(190) xor d(189) xor d(188) xor d(187) xor d(185) xor d(183) xor d(180) xor d(179) xor d(169) xor d(168) xor d(167) xor d(166) xor d(164) xor d(163) xor d(159) xor d(158) xor d(155) xor d(153) xor d(152) xor d(148) xor d(146) xor d(141) xor d(140) xor d(134) xor d(133) xor d(132) xor d(131) xor d(129) xor d(125) xor d(124) xor d(123) xor d(122) xor d(120) xor d(116) xor d(115) xor d(114) xor d(113) xor d(111) xor d(110) xor d(108) xor d(107) xor d(103) xor d(101) xor d(100) xor d(98) xor d(96) xor d(95) xor d(94) xor d(93) xor d(92) xor d(91) xor d(84) xor d(82) xor d(81) xor d(80) xor d(79) xor d(78) xor d(76) xor d(70) xor d(69) xor d(65) xor d(64) xor d(63) xor d(62) xor d(60) xor d(58) xor d(57) xor d(55) xor d(52) xor d(51) xor d(50) xor d(47) xor d(45) xor d(44) xor d(42) xor d(41) xor d(34) xor d(31) xor d(29) xor d(28) xor d(27) xor d(26) xor d(25) xor d(23) xor d(22) xor d(21) xor d(13) xor d(9) xor d(7) xor d(6) xor d(3) xor c(0) xor c(3) xor c(5) xor c(6) xor c(7) xor c(8) xor c(9) xor c(10) xor c(11) xor c(12) xor c(17) xor c(18) xor c(19) xor c(23) xor c(24) xor c(25) xor c(27) xor c(28) xor c(29) xor c(31);
    newcrc(30) := d(510) xor d(509) xor d(508) xor d(506) xor d(505) xor d(504) xor d(500) xor d(499) xor d(498) xor d(493) xor d(492) xor d(491) xor d(490) xor d(489) xor d(488) xor d(487) xor d(486) xor d(484) xor d(481) xor d(480) xor d(479) xor d(478) xor d(477) xor d(475) xor d(474) xor d(470) xor d(468) xor d(466) xor d(463) xor d(462) xor d(460) xor d(459) xor d(456) xor d(450) xor d(448) xor d(447) xor d(446) xor d(442) xor d(435) xor d(434) xor d(432) xor d(431) xor d(422) xor d(420) xor d(417) xor d(416) xor d(414) xor d(412) xor d(410) xor d(407) xor d(406) xor d(405) xor d(403) xor d(402) xor d(398) xor d(397) xor d(396) xor d(394) xor d(391) xor d(390) xor d(389) xor d(388) xor d(386) xor d(385) xor d(384) xor d(379) xor d(376) xor d(374) xor d(372) xor d(370) xor d(367) xor d(366) xor d(364) xor d(361) xor d(360) xor d(357) xor d(356) xor d(355) xor d(351) xor d(347) xor d(346) xor d(345) xor d(343) xor d(342) xor d(340) xor d(339) xor d(337) xor d(336) xor d(335) xor d(333) xor d(332) xor d(331) xor d(326) xor d(325) xor d(320) xor d(319) xor d(318) xor d(317) xor d(316) xor d(315) xor d(313) xor d(310) xor d(308) xor d(307) xor d(303) xor d(301) xor d(300) xor d(298) xor d(297) xor d(296) xor d(295) xor d(294) xor d(293) xor d(292) xor d(290) xor d(288) xor d(286) xor d(285) xor d(284) xor d(281) xor d(277) xor d(275) xor d(274) xor d(272) xor d(271) xor d(267) xor d(266) xor d(263) xor d(262) xor d(259) xor d(257) xor d(255) xor d(253) xor d(250) xor d(246) xor d(241) xor d(235) xor d(232) xor d(228) xor d(226) xor d(225) xor d(224) xor d(222) xor d(214) xor d(212) xor d(210) xor d(208) xor d(207) xor d(206) xor d(205) xor d(201) xor d(200) xor d(199) xor d(197) xor d(196) xor d(195) xor d(192) xor d(191) xor d(190) xor d(189) xor d(188) xor d(186) xor d(184) xor d(181) xor d(180) xor d(170) xor d(169) xor d(168) xor d(167) xor d(165) xor d(164) xor d(160) xor d(159) xor d(156) xor d(154) xor d(153) xor d(149) xor d(147) xor d(142) xor d(141) xor d(135) xor d(134) xor d(133) xor d(132) xor d(130) xor d(126) xor d(125) xor d(124) xor d(123) xor d(121) xor d(117) xor d(116) xor d(115) xor d(114) xor d(112) xor d(111) xor d(109) xor d(108) xor d(104) xor d(102) xor d(101) xor d(99) xor d(97) xor d(96) xor d(95) xor d(94) xor d(93) xor d(92) xor d(85) xor d(83) xor d(82) xor d(81) xor d(80) xor d(79) xor d(77) xor d(71) xor d(70) xor d(66) xor d(65) xor d(64) xor d(63) xor d(61) xor d(59) xor d(58) xor d(56) xor d(53) xor d(52) xor d(51) xor d(48) xor d(46) xor d(45) xor d(43) xor d(42) xor d(35) xor d(32) xor d(30) xor d(29) xor d(28) xor d(27) xor d(26) xor d(24) xor d(23) xor d(22) xor d(14) xor d(10) xor d(8) xor d(7) xor d(4) xor c(0) xor c(1) xor c(4) xor c(6) xor c(7) xor c(8) xor c(9) xor c(10) xor c(11) xor c(12) xor c(13) xor c(18) xor c(19) xor c(20) xor c(24) xor c(25) xor c(26) xor c(28) xor c(29) xor c(30);
    newcrc(31) := d(511) xor d(510) xor d(509) xor d(507) xor d(506) xor d(505) xor d(501) xor d(500) xor d(499) xor d(494) xor d(493) xor d(492) xor d(491) xor d(490) xor d(489) xor d(488) xor d(487) xor d(485) xor d(482) xor d(481) xor d(480) xor d(479) xor d(478) xor d(476) xor d(475) xor d(471) xor d(469) xor d(467) xor d(464) xor d(463) xor d(461) xor d(460) xor d(457) xor d(451) xor d(449) xor d(448) xor d(447) xor d(443) xor d(436) xor d(435) xor d(433) xor d(432) xor d(423) xor d(421) xor d(418) xor d(417) xor d(415) xor d(413) xor d(411) xor d(408) xor d(407) xor d(406) xor d(404) xor d(403) xor d(399) xor d(398) xor d(397) xor d(395) xor d(392) xor d(391) xor d(390) xor d(389) xor d(387) xor d(386) xor d(385) xor d(380) xor d(377) xor d(375) xor d(373) xor d(371) xor d(368) xor d(367) xor d(365) xor d(362) xor d(361) xor d(358) xor d(357) xor d(356) xor d(352) xor d(348) xor d(347) xor d(346) xor d(344) xor d(343) xor d(341) xor d(340) xor d(338) xor d(337) xor d(336) xor d(334) xor d(333) xor d(332) xor d(327) xor d(326) xor d(321) xor d(320) xor d(319) xor d(318) xor d(317) xor d(316) xor d(314) xor d(311) xor d(309) xor d(308) xor d(304) xor d(302) xor d(301) xor d(299) xor d(298) xor d(297) xor d(296) xor d(295) xor d(294) xor d(293) xor d(291) xor d(289) xor d(287) xor d(286) xor d(285) xor d(282) xor d(278) xor d(276) xor d(275) xor d(273) xor d(272) xor d(268) xor d(267) xor d(264) xor d(263) xor d(260) xor d(258) xor d(256) xor d(254) xor d(251) xor d(247) xor d(242) xor d(236) xor d(233) xor d(229) xor d(227) xor d(226) xor d(225) xor d(223) xor d(215) xor d(213) xor d(211) xor d(209) xor d(208) xor d(207) xor d(206) xor d(202) xor d(201) xor d(200) xor d(198) xor d(197) xor d(196) xor d(193) xor d(192) xor d(191) xor d(190) xor d(189) xor d(187) xor d(185) xor d(182) xor d(181) xor d(171) xor d(170) xor d(169) xor d(168) xor d(166) xor d(165) xor d(161) xor d(160) xor d(157) xor d(155) xor d(154) xor d(150) xor d(148) xor d(143) xor d(142) xor d(136) xor d(135) xor d(134) xor d(133) xor d(131) xor d(127) xor d(126) xor d(125) xor d(124) xor d(122) xor d(118) xor d(117) xor d(116) xor d(115) xor d(113) xor d(112) xor d(110) xor d(109) xor d(105) xor d(103) xor d(102) xor d(100) xor d(98) xor d(97) xor d(96) xor d(95) xor d(94) xor d(93) xor d(86) xor d(84) xor d(83) xor d(82) xor d(81) xor d(80) xor d(78) xor d(72) xor d(71) xor d(67) xor d(66) xor d(65) xor d(64) xor d(62) xor d(60) xor d(59) xor d(57) xor d(54) xor d(53) xor d(52) xor d(49) xor d(47) xor d(46) xor d(44) xor d(43) xor d(36) xor d(33) xor d(31) xor d(30) xor d(29) xor d(28) xor d(27) xor d(25) xor d(24) xor d(23) xor d(15) xor d(11) xor d(9) xor d(8) xor d(5) xor c(0) xor c(1) xor c(2) xor c(5) xor c(7) xor c(8) xor c(9) xor c(10) xor c(11) xor c(12) xor c(13) xor c(14) xor c(19) xor c(20) xor c(21) xor c(25) xor c(26) xor c(27) xor c(29) xor c(30) xor c(31);
    return newcrc;
  end nextCRC32_D512;

end PCK_CRC32_D512;
