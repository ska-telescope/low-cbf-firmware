--
-- FB_top.vhd
-- Author : David Humphrey (dave.humphrey@csiro.au)
-- Description
--  Top level for the perentie filterbanks. Includes :
--   - Correlator filterbank - 4096 point FFT, 12 tap FIR filter, 4 streams simultaneously.
--   - PSS filterbank - 64 point FFT, 12 tap FIR filter, 6 streams simultaneously.
--   - PST filterbank - 256 point FFT, 12 tap FIR filter, oversampled by 4/3, 6 streams simultaneously.
--   - MACE interface, which is just to allow reading/writing of the filter taps in the filterbanks.
--     *** WARNING *** MACE slave is manually written. MACE slave module is NOT auto-generated by ARGS. 
--     Changing the yaml file will not change the actual registers.
--     This is to allow the memories to reside in the filters, rather than being pulled out and put into 
--     ARGs. 
--
----------------------------------------------------------------------------------------------------------
library IEEE, axi4_lib, ctc_lib, common_lib, filterbanks_lib;
use ctc_lib.ctc_pkg.all;
use common_lib.common_pkg.all;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use axi4_lib.axi4_lite_pkg.ALL;
use axi4_lib.axi4_full_pkg.ALL;
--USE filterbanks_lib.filterbanks_reg_pkg.ALL;

entity FB_Top is
    generic(
        USE_CORRELATOR_FB : boolean := true;
        USE_PSS_FB : boolean := true;
        USE_PST_FB : boolean := true
    );
    port(
        -- clock, target is 400 MHz
        i_data_clk       : in std_logic;
        i_data_rst       : in std_logic;
        -- AXI slave interface, 64k word block of space with the fir filter coefficients.
        i_MACE_clk  : in std_logic;
        i_MACE_rst  : in std_logic;
        i_axi_mosi  : in  t_axi4_full_mosi;
        o_axi_miso  : out t_axi4_full_miso;
        -----------------------------------------
        -- Correlator filterbank input.
        i_CorSOF         : in std_logic;                            -- start of frame.
        i_CorHeader      : in t_ctc_output_header_a(1 downto 0);    -- meta data belonging to the data coming out
        i_CorHeaderValid : in std_logic;                            -- new meta data (every output packet, aka 4096 cycles) 
        i_CorData        : in t_ctc_output_data_a(1 downto 0);      -- the actual output data
        i_CorDataValid   : in std_logic;
        -- Correlator Filterbank output
        o_CorHeader      : out t_ctc_output_header_a(1 downto 0);    -- meta data belonging to the data coming out
        o_CorHeaderValid : out std_logic;                            -- new meta data (every output packet, aka 4096 cycles) 
        o_CorData        : out t_ctc_output_data_a(1 downto 0);      -- the actual output data
        o_CorDataValid   : out std_logic;
        -----------------------------------------
        -- PSS and PST Data input, common valid signal, expects packets of 64 samples. 
        -- Requires at least 2 clocks idle time between packets.
        -- Due to oversampling, also requires on average 86 clocks between packets - specifically, no more than 3 packets in 258 clocks.
        i_PSSPSTSOF         : in std_logic; 
        i_PSSPSTHeader      : in t_ctc_output_header_a(2 downto 0);
        i_PSSPSTHeaderValid : in std_logic;
        i_PSSPSTData        : in t_ctc_output_data_a(2 downto 0);
        i_PSSPSTDataValid   : in std_logic;
        -- PSS filterbank data Output
        o_PSSHeader      : out t_ctc_output_header_a(2 downto 0);
        o_PSSHeaderValid : out std_logic;
        o_PSSData        : out t_ctc_output_data_a(2 downto 0);
        o_PSSDataValid   : out std_logic;
        -- PST filterbank data output
        o_PSTHeader      : out t_ctc_output_header_a(2 downto 0);
        o_PSTHeaderValid : out std_logic;
        o_PSTData        : out t_ctc_output_data_a(2 downto 0);
        o_PSTDataValid   : out std_logic
    );
end FB_Top;

architecture Behavioral of FB_Top is
    
    signal firtap_addr : std_logic_vector(15 downto 0);
    signal firtap_clk : std_logic;
    signal cor_we : std_logic;
    signal PSS_we : std_logic;
    signal PST_we : std_logic;
    signal corFirRd_data : std_logic_vector(17 downto 0);
    signal PSTfirRd_data : std_logic_vector(17 downto 0);
    signal PSSfirRd_data : std_logic_vector(17 downto 0);
    signal firtap_wr_data : std_logic_vector(17 downto 0);
    
    signal CorDin0, CorDin1, CorDin2, CorDin3 : t_slv_8_arr(1 downto 0);
    signal CorMetaIn, CorMetaOut : std_logic_vector(209 downto 0);
    signal CorDout0, CorDout1, CorDout2, CorDout3 : t_slv_16_arr(1 downto 0);
    signal CorValidOut, CorValidOutDel : std_logic;
    
    signal PSSPSTDin0, PSSPSTDin1, PSSPSTDin2, PSSPSTDin3, PSSPSTDin4, PSSPSTDin5 : t_slv_8_arr(1 downto 0);
    signal PSSPSTMetaIn, PSSMetaOut, PSTMetaOut : std_logic_vector(314 downto 0);
    signal PSTDout0, PSTDout1, PSTDout2, PSTDout3, PSTDout4, PSTDout5 : t_slv_16_arr(1 downto 0);
    signal PSSDout0, PSSDout1, PSSDout2, PSSDout3, PSSDout4, PSSDout5 : t_slv_16_arr(1 downto 0);
    signal PSSValidOut, PSTValidOut, PSSValidOutDel, PSTValidOutDel : std_logic;
    
begin
    
    -----------------------------------------------------------------------------------
    -- Correlator Filterbank
    --
    -- Note : 
    --    type t_ctc_output_header is record
    --        timestamp         : std_logic_vector(42 downto 0);
    --        coarse_delay      : std_logic_vector(11 downto 0);
    --        virtual_channel   : std_logic_vector(8 downto 0);
    --        station_id        : std_logic_vector(8 downto 0);
    --        hpol_phase_shift  : std_logic_vector(15 downto 0);  
    --        vpol_phase_shift  : std_logic_vector(15 downto 0);  
    --    end record;
    
    CorDin0(0) <= i_CorData(0).data.vpol.re;
    CorDin0(1) <= i_CorData(0).data.vpol.im;
    CorDin1(0) <= i_CorData(0).data.hpol.re;
    CorDin1(1) <= i_CorData(0).data.hpol.im;
    CorDin2(0) <= i_CorData(1).data.vpol.re;
    CorDin2(1) <= i_CorData(1).data.vpol.im;
    CorDin3(0) <= i_CorData(1).data.hpol.re;
    CorDin3(1) <= i_CorData(1).data.hpol.im;
    CorMetaIn(42 downto 0) <= i_CorHeader(0).timestamp; -- 43 bits
    CorMetaIn(54 downto 43) <= i_CorHeader(0).coarse_delay; -- 12 bits
    CorMetaIn(63 downto 55) <= i_CorHeader(0).virtual_channel; -- 9 bits
    CorMetaIn(72 downto 64) <= i_CorHeader(0).station_id; -- 9 bits 
    CorMetaIn(88 downto 73) <= i_CorHeader(0).hpol_phase_shift; -- 16 bits
    CorMetaIn(104 downto 89) <= i_CorHeader(0).vpol_phase_shift; -- 16 bits
    CorMetaIn(42+105 downto 0+105) <= i_CorHeader(1).timestamp; -- 43 bits
    CorMetaIn(54+105 downto 43+105) <= i_CorHeader(1).coarse_delay; -- 12 bits
    CorMetaIn(63+105 downto 55+105) <= i_CorHeader(1).virtual_channel; -- 9 bits
    CorMetaIn(72+105 downto 64+105) <= i_CorHeader(1).station_id; -- 9 bits 
    CorMetaIn(88+105 downto 73+105) <= i_CorHeader(1).hpol_phase_shift; -- 16 bits
    CorMetaIn(104+105 downto 89+105) <= i_CorHeader(1).vpol_phase_shift; -- 16 bits
    
    corfbi : entity filterbanks_lib.correlatorFBTop25
    generic map (
        METABITS => 210,    --  integer := 64; -- Width in bits of the meta_i and meta_o ports.
        FRAMESTODROP => 11  --  integer := 11  -- Number of output frames to drop after a reset (to account for initialisation of the filterbank)
    )
    port map(
        -- clock, target is 380 MHz
        clk => i_data_clk,  -- in std_logic;
        rst => i_corSOF,    -- in std_logic;
        -- Data input, common valid signal, expects packets of 4096 samples. Requires at least 2 clocks idle time between packets.
        data0_i => CorDin0,        -- in t_slv_8_arr(1:0); 4 Inputs, each complex data, 8 bit real, 8 bit imaginary.
        data1_i => CorDin1,        -- in t_slv_8_arr(1:0);
        data2_i => CorDin2,        -- in t_slv_8_arr(1:0);
        data3_i => CorDin2,        -- in t_slv_8_arr(1:0);
        meta_i  => CorMetaIn,        -- in ((METABITS-1) downto 0);
        valid_i => i_CorDataValid, -- in std_logic;
        -- Data out; bursts of 3456 clocks for each channel.
        data0_o => CorDout0,    -- out t_slv_16_arr(1 downto 0);   -- 4 outputs, real and imaginary parts in (0) and (1) respectively;
        data1_o => CorDout1,    -- out t_slv_16_arr(1 downto 0);
        data2_o => CorDout2,    -- out t_slv_16_arr(1 downto 0);
        data3_o => CorDout3,    -- out t_slv_16_arr(1 downto 0);
        meta_o  => CorMetaOut,  -- out std_logic_vector((METABITS-1) downto 0);
        valid_o => CorValidOut, -- out std_logic;
        -- Writing FIR Taps
        FIRTapData_i => firtap_wr_data, --: in std_logic_vector(17 downto 0);  -- For register writes of the filtertaps.
        FIRTapData_o => corFirRd_data, -- : out std_logic_vector(17 downto 0); -- For register reads of the filtertaps. 3 cycle latency from FIRTapAddr_i
        FIRTapAddr_i => firtap_addr(15 downto 0), --: in std_logic_vector(15 downto 0);  -- 4096 * 12 filter taps = 49152 total.
        FIRTapWE_i   => cor_we, -- : in std_logic;
        FIRTapClk    => firtap_clk --: in std_logic
    );

    -- Just use the low 8 bits; need to replace this with the RFI module.
    o_CorData(0).data.vpol.re <= CorDout0(0)(7 downto 0);
    o_CorData(0).data.vpol.im <= CorDout0(1)(7 downto 0);
    o_CorData(0).data.hpol.re <= CorDout1(0)(7 downto 0);
    o_CorData(0).data.hpol.im <= CorDout1(1)(7 downto 0);
    o_CorData(1).data.vpol.re <= CorDout2(0)(7 downto 0);
    o_CorData(1).data.vpol.im <= CorDout2(1)(7 downto 0);
    o_CorData(1).data.hpol.re <= CorDout3(0)(7 downto 0);
    o_CorData(1).data.hpol.im <= CorDout3(1)(7 downto 0);
    o_CorDataValid <= CorValidOut;
    
    o_CorHeader(0).timestamp        <= CorMetaOut(42 downto 0);
    o_CorHeader(0).coarse_delay     <= CorMetaOut(54 downto 43);
    o_CorHeader(0).virtual_channel  <= CorMetaOut(63 downto 55);
    o_CorHeader(0).station_id       <= CorMetaOut(72 downto 64); 
    o_CorHeader(0).hpol_phase_shift <= CorMetaOut(88 downto 73);
    o_CorHeader(0).vpol_phase_shift <= CorMetaOut(104 downto 89);
    o_CorHeader(1).timestamp        <= CorMetaOut(42+105 downto 0+105);
    o_CorHeader(1).coarse_delay     <= CorMetaOut(54+105 downto 43+105);
    o_CorHeader(1).virtual_channel  <= CorMetaOut(63+105 downto 55+105);
    o_CorHeader(1).station_id       <= CorMetaOut(72+105 downto 64+105); 
    o_CorHeader(1).hpol_phase_shift <= CorMetaOut(88+105 downto 73+105);
    o_CorHeader(1).vpol_phase_shift <= CorMetaOut(104+105 downto 89+105);
    o_CorHeaderValid <= CorValidOut and (not CorValidOutDel);
    
    process(i_data_clk)
    begin
        if rising_edge(i_data_clk) then
            CorValidOutDel <= CorValidOut;
        end if;
    end process;
    
    -----------------------------------------------------------------------------------
    -- PST Filterbank
    PSSPSTDin0(0) <= i_PSSPSTData(0).data.vpol.re;
    PSSPSTDin0(1) <= i_PSSPSTData(0).data.vpol.im;
    PSSPSTDin1(0) <= i_PSSPSTData(0).data.hpol.re;
    PSSPSTDin1(1) <= i_PSSPSTData(0).data.hpol.im;
    PSSPSTDin2(0) <= i_PSSPSTData(1).data.vpol.re;
    PSSPSTDin2(1) <= i_PSSPSTData(1).data.vpol.im;
    PSSPSTDin3(0) <= i_PSSPSTData(1).data.hpol.re;
    PSSPSTDin3(1) <= i_PSSPSTData(1).data.hpol.im;
    PSSPSTDin4(0) <= i_PSSPSTData(2).data.vpol.re;
    PSSPSTDin4(1) <= i_PSSPSTData(2).data.vpol.im;
    PSSPSTDin5(0) <= i_PSSPSTData(2).data.hpol.re;
    PSSPSTDin5(1) <= i_PSSPSTData(2).data.hpol.im;
    
    PSSPSTMetaIn(42 downto 0) <= i_PSSPSTHeader(0).timestamp; -- 43 bits
    PSSPSTMetaIn(54 downto 43) <= i_PSSPSTHeader(0).coarse_delay; -- 12 bits
    PSSPSTMetaIn(63 downto 55) <= i_PSSPSTHeader(0).virtual_channel; -- 9 bits
    PSSPSTMetaIn(72 downto 64) <= i_PSSPSTHeader(0).station_id; -- 9 bits 
    PSSPSTMetaIn(88 downto 73) <= i_PSSPSTHeader(0).hpol_phase_shift; -- 16 bits
    PSSPSTMetaIn(104 downto 89) <= i_PSSPSTHeader(0).vpol_phase_shift; -- 16 bits
    PSSPSTMetaIn(42+105 downto 0+105) <= i_PSSPSTHeader(1).timestamp; -- 43 bits
    PSSPSTMetaIn(54+105 downto 43+105) <= i_PSSPSTHeader(1).coarse_delay; -- 12 bits
    PSSPSTMetaIn(63+105 downto 55+105) <= i_PSSPSTHeader(1).virtual_channel; -- 9 bits
    PSSPSTMetaIn(72+105 downto 64+105) <= i_PSSPSTHeader(1).station_id; -- 9 bits 
    PSSPSTMetaIn(88+105 downto 73+105) <= i_PSSPSTHeader(1).hpol_phase_shift; -- 16 bits
    PSSPSTMetaIn(104+105 downto 89+105) <= i_PSSPSTHeader(1).vpol_phase_shift; -- 16 bits
    PSSPSTMetaIn(42+210 downto 0+210) <= i_PSSPSTHeader(2).timestamp; -- 43 bits
    PSSPSTMetaIn(54+210 downto 43+210) <= i_PSSPSTHeader(2).coarse_delay; -- 12 bits
    PSSPSTMetaIn(63+210 downto 55+210) <= i_PSSPSTHeader(2).virtual_channel; -- 9 bits
    PSSPSTMetaIn(72+210 downto 64+210) <= i_PSSPSTHeader(2).station_id; -- 9 bits 
    PSSPSTMetaIn(88+210 downto 73+210) <= i_PSSPSTHeader(2).hpol_phase_shift; -- 16 bits
    PSSPSTMetaIn(104+210 downto 89+210) <= i_PSSPSTHeader(2).vpol_phase_shift; -- 16 bits    
    
    
    pstfbi : entity filterbanks_lib.PSTFBTop
    generic map(
        METABITS => 315,    -- Width in bits of the meta_i and meta_o ports.
        FRAMESTODROP => 11  -- Number of output frames to drop after a reset (to account for initialisation of the filterbank)
    )
    port map (
        -- processing clock
        clk         => i_data_clk,
        rst         => i_PSSPSTSOF,
        FIRTapUse_i => '0', --in std_logic; FIR Taps are double buffered, choose which set of TAPs to use.
        -- Data input, common valid signal, expects packets of 64 samples. 
        -- Requires at least 2 clocks idle time between packets.
        -- Due to oversampling, also requires on average 86 clocks between packets - specifically, no more than 3 packets in 258 clocks. 
        data0_i => PSSPSTDin0, -- in t_slv_8_arr(1 downto 0);  -- 6 Inputs, each complex data, 8 bit real, 8 bit imaginary.
        data1_i => PSSPSTDin1, -- in t_slv_8_arr(1 downto 0);
        data2_i => PSSPSTDin2, -- in t_slv_8_arr(1 downto 0);
        data3_i => PSSPSTDin3, -- in t_slv_8_arr(1 downto 0);
        data4_i => PSSPSTDin4, -- in t_slv_8_arr(1 downto 0);
        data5_i => PSSPSTDin5, -- in t_slv_8_arr(1 downto 0);
        meta_i  => PSSPSTMetaIn, -- in std_logic_vector((METABITS-1) downto 0);  -- Sampled on the first cycle of every third packet of valid_i. 
        valid_i => i_PSSPSTDataValid, -- in std_logic;
        -- Data out; bursts of 216 clocks for each channel.
        data0_o => PSTDout0,    -- out t_slv_16_arr(1 downto 0);   -- 6 outputs, real and imaginary parts in (0) and (1) respectively;
        data1_o => PSTDout1,    -- out t_slv_16_arr(1 downto 0);
        data2_o => PSTDout2,    -- out t_slv_16_arr(1 downto 0);
        data3_o => PSTDout3,    -- out t_slv_16_arr(1 downto 0);
        data4_o => PSTDout4,    -- out t_slv_16_arr(1 downto 0);
        data5_o => PSTDout5,    -- out t_slv_16_arr(1 downto 0);
        meta_o  => PSTMetaOut,  -- out std_logic_vector((METABITS-1) downto 0);
        valid_o => PSTValidOut, -- out std_logic;
        -- Writing FIR Taps
        FIRTapData_i   => firtap_wr_data, --: in std_logic_vector(17 downto 0);  -- For register writes of the filtertaps.
        FIRTapData_o   => PSTfirRd_data, -- : out std_logic_vector(17 downto 0); -- For register reads of the filtertaps. 3 cycle latency from FIRTapAddr_i
        FIRTapAddr_i   => firtap_addr(11 downto 0), --: in std_logic_vector(11 downto 0);   -- 256 * 12 filter taps = 3072 total.
        FIRTapWE_i     => PST_we, -- : in std_logic;
        FIRTapClk      => firtap_clk, --: in std_logic;
        FIRTapSelect_i => '0' -- : in std_logic  -- FIR Taps are double buffered; This selects the buffer to access for registers. Choose which buffer to use with FIRTapUse_i
    );

    -- Just use the low 8 bits; need to replace this with the RFI module.
    o_PSTData(0).data.vpol.re <= PSTDout0(0)(7 downto 0);
    o_PSTData(0).data.vpol.im <= PSTDout0(1)(7 downto 0);
    o_PSTData(0).data.hpol.re <= PSTDout1(0)(7 downto 0);
    o_PSTData(0).data.hpol.im <= PSTDout1(1)(7 downto 0);
    o_PSTData(1).data.vpol.re <= PSTDout2(0)(7 downto 0);
    o_PSTData(1).data.vpol.im <= PSTDout2(1)(7 downto 0);
    o_PSTData(1).data.hpol.re <= PSTDout3(0)(7 downto 0);
    o_PSTData(1).data.hpol.im <= PSTDout3(1)(7 downto 0);
    o_PSTData(2).data.vpol.re <= PSTDout4(0)(7 downto 0);
    o_PSTData(2).data.vpol.im <= PSTDout4(1)(7 downto 0);
    o_PSTData(2).data.hpol.re <= PSTDout5(0)(7 downto 0);
    o_PSTData(2).data.hpol.im <= PSTDout5(1)(7 downto 0);
    o_PSTDataValid <= PSTValidOut;
    
    o_PSTHeader(0).timestamp        <= PSTMetaOut(42 downto 0);
    o_PSTHeader(0).coarse_delay     <= PSTMetaOut(54 downto 43);
    o_PSTHeader(0).virtual_channel  <= PSTMetaOut(63 downto 55);
    o_PSTHeader(0).station_id       <= PSTMetaOut(72 downto 64); 
    o_PSTHeader(0).hpol_phase_shift <= PSTMetaOut(88 downto 73);
    o_PSTHeader(0).vpol_phase_shift <= PSTMetaOut(104 downto 89);
    o_PSTHeader(1).timestamp        <= PSTMetaOut(42+105 downto 0+105);
    o_PSTHeader(1).coarse_delay     <= PSTMetaOut(54+105 downto 43+105);
    o_PSTHeader(1).virtual_channel  <= PSTMetaOut(63+105 downto 55+105);
    o_PSTHeader(1).station_id       <= PSTMetaOut(72+105 downto 64+105); 
    o_PSTHeader(1).hpol_phase_shift <= PSTMetaOut(88+105 downto 73+105);
    o_PSTHeader(1).vpol_phase_shift <= PSTMetaOut(104+105 downto 89+105);
    o_PSTHeader(2).timestamp        <= PSTMetaOut(42+210 downto 0+210);
    o_PSTHeader(2).coarse_delay     <= PSTMetaOut(54+210 downto 43+210);
    o_PSTHeader(2).virtual_channel  <= PSTMetaOut(63+210 downto 55+210);
    o_PSTHeader(2).station_id       <= PSTMetaOut(72+210 downto 64+210); 
    o_PSTHeader(2).hpol_phase_shift <= PSTMetaOut(88+210 downto 73+210);
    o_PSTHeader(2).vpol_phase_shift <= PSTMetaOut(104+210 downto 89+210);
    
    o_PSTHeaderValid <= PSTValidOut and (not PSTValidOutDel);
    
    process(i_data_clk)
    begin
        if rising_edge(i_data_clk) then
            PSTValidOutDel <= PSTValidOut;
        end if;
    end process;

    
    pssfbi : entity filterbanks_lib.PSSFBTop
    port map(
        -- processing clock
        clk         => i_data_clk,
        rst         => i_PSSPSTSOF,
        FIRTapUse_i => '0', -- : in std_logic;   -- FIR Taps are double buffered, choose which set of TAPs to use.
        -- Data input, common valid signal, expects packets of 64 samples. Requires at least 2 clocks idle time between packets.
        data0_i => PSSPSTDin0, -- in t_slv_8_arr(1 downto 0);  -- 6 Inputs, each complex data, 8 bit real, 8 bit imaginary.
        data1_i => PSSPSTDin1, -- in t_slv_8_arr(1 downto 0);
        data2_i => PSSPSTDin2, -- in t_slv_8_arr(1 downto 0);
        data3_i => PSSPSTDin3, -- in t_slv_8_arr(1 downto 0);
        data4_i => PSSPSTDin4, -- in t_slv_8_arr(1 downto 0);
        data5_i => PSSPSTDin5, -- in t_slv_8_arr(1 downto 0);
        valid_i => i_PSSPSTDataValid, -- in std_logic;
        -- Data out; bursts of 54 clocks for each channel.
        data0_o => PSSDout0,    -- out t_slv_16_arr(1 downto 0);   -- 6 outputs, real and imaginary parts in (0) and (1) respectively;
        data1_o => PSSDout1,    -- out t_slv_16_arr(1 downto 0);
        data2_o => PSSDout2,    -- out t_slv_16_arr(1 downto 0);
        data3_o => PSSDout3,    -- out t_slv_16_arr(1 downto 0);
        data4_o => PSSDout4,    -- out t_slv_16_arr(1 downto 0);
        data5_o => PSSDout5,    -- out t_slv_16_arr(1 downto 0);
        valid_o => PSSValidOut,  -- out std_logic;
        -- Writing FIR Taps
        FIRTapData_i   => firtap_wr_data, --: in std_logic_vector(17 downto 0);  -- For register writes of the filtertaps.
        FIRTapData_o   => PSSfirRd_data, --: out std_logic_vector(17 downto 0); -- For register reads of the filtertaps. 3 cycle latency from FIRTapAddr_i
        FIRTapAddr_i   => firtap_addr(9 downto 0), -- : in std_logic_vector(9 downto 0);   -- 64 * 12 filter taps = 768 total.
        FIRTapWE_i     => PSS_we, -- : in std_logic;
        FIRTapClk      => firtap_clk, --  in std_logic;
        FIRTapSelect_i => '0' -- : in std_logic  -- FIR Taps are double buffered; This selects the buffer to access for registers. Choose which buffer to use with FIRTapUse_i
    );

    -- Just use the low 8 bits; need to replace this with the RFI module.
    o_PSSData(0).data.vpol.re <= PSSDout0(0)(7 downto 0);
    o_PSSData(0).data.vpol.im <= PSSDout0(1)(7 downto 0);
    o_PSSData(0).data.hpol.re <= PSSDout1(0)(7 downto 0);
    o_PSSData(0).data.hpol.im <= PSSDout1(1)(7 downto 0);
    o_PSSData(1).data.vpol.re <= PSSDout2(0)(7 downto 0);
    o_PSSData(1).data.vpol.im <= PSSDout2(1)(7 downto 0);
    o_PSSData(1).data.hpol.re <= PSSDout3(0)(7 downto 0);
    o_PSSData(1).data.hpol.im <= PSSDout3(1)(7 downto 0);
    o_PSSData(2).data.vpol.re <= PSSDout4(0)(7 downto 0);
    o_PSSData(2).data.vpol.im <= PSSDout4(1)(7 downto 0);
    o_PSSData(2).data.hpol.re <= PSSDout5(0)(7 downto 0);
    o_PSSData(2).data.hpol.im <= PSSDout5(1)(7 downto 0);
    o_PSSDataValid <= PSSValidOut;
    
    -- To be fixed...
    o_PSSHeader(0).timestamp        <= (others => '0');
    o_PSSHeader(0).coarse_delay     <= (others => '0');
    o_PSSHeader(0).virtual_channel  <= (others => '0');
    o_PSSHeader(0).station_id       <= (others => '0');
    o_PSSHeader(0).hpol_phase_shift <= (others => '0');
    o_PSSHeader(0).vpol_phase_shift <= (others => '0');
    o_PSSHeader(1).timestamp        <= (others => '0');
    o_PSSHeader(1).coarse_delay     <= (others => '0');
    o_PSSHeader(1).virtual_channel  <= (others => '0');
    o_PSSHeader(1).station_id       <= (others => '0');
    o_PSSHeader(1).hpol_phase_shift <= (others => '0');
    o_PSSHeader(1).vpol_phase_shift <= (others => '0');
    o_PSSHeader(2).timestamp        <= (others => '0');
    o_PSSHeader(2).coarse_delay     <= (others => '0');
    o_PSSHeader(2).virtual_channel  <= (others => '0');
    o_PSSHeader(2).station_id       <= (others => '0');
    o_PSSHeader(2).hpol_phase_shift <= (others => '0');
    o_PSSHeader(2).vpol_phase_shift <= (others => '0'); 
    
    o_PSSHeaderValid <= PSSValidOut and (not PSSValidOutDel);
    
    process(i_data_clk)
    begin
        if rising_edge(i_data_clk) then
            PSSValidOutDel <= PSSValidOut;
        end if;
    end process;
    
    ---------------------------------------------------------------
    -- Programming the FIR taps in the filters
    
    mmfirtapsi : entity filterbanks_lib.filterbanks_firtaps_ram
    port map (
        -- full AXI bus
        CLK_A      => i_MACE_clk, -- IN  STD_LOGIC;
        RST_A      => i_MACE_rst, -- IN  STD_LOGIC;
        MM_IN      => i_axi_mosi, -- IN  t_axi4_full_mosi;
        MM_OUT     => o_axi_miso, -- OUT t_axi4_full_miso;
        -- Interface to the memories. Should be a 3 cycle latency for reads
        -- Note - two extra cycles of latency added in this file, so axi interface is configured for 5 cycle read latency.
        -- Common memory interface signals
        mem_clk    => firtap_clk,  -- out std_logic;
        mem_rst    => open,        -- out std_logic;
        mem_addr   => firtap_addr, -- out std_logic_vector(15 downto 0);
        mem_wr_data => firtap_wr_data, --  out std_logic_vector(17 downto 0);
        -- Correlator - address 0 to 49151 (0x0 to 0xC000)
        o_cor_we     => cor_we, -- : out std_logic;
        i_cor_rd_data => corFirRd_data, -- : in std_logic_vector(17 downto 0);
        -- PST - 3072 words, address 49152 to 52223 (0xC000 to 0xCBFF)
        o_PST_we => PST_we, -- : out std_logic;
        i_PST_rd_data => PSTfirRd_data, -- : in std_logic_vector(17 downto 0);
        -- PSS - 768 words, Address 53248 to 54015 (0xD000 to 0xD2FF)
        o_PSS_we  => PSS_we, -- : out std_logic;
        i_PSS_rd_data => PSSfirRd_data -- : in std_logic_vector(17 downto 0)
    ); 
    
    
end Behavioral;