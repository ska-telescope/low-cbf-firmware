--------------------------------------------------------------------------------
-- Copyright (C) 1999-2008 Easics NV.
-- This source file may be used and distributed without restriction
-- provided that this copyright statement is not removed from the file
-- and that any derivative work contains the original copyright notice
-- and the associated disclaimer.
--
-- THIS SOURCE FILE IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS
-- OR IMPLIED WARRANTIES, INCLUDING, WITHOUT LIMITATION, THE IMPLIED
-- WARRANTIES OF MERCHANTIBILITY AND FITNESS FOR A PARTICULAR PURPOSE.
--
-- Purpose : synthesizable CRC function
--   * polynomial: (0 1 2 4 5 7 8 10 11 12 16 22 23 26 32)
--   * data width: 1024
--
-- Info : tools@easics.be
--        http://www.easics.com
--------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

package PCK_CRC32_D1024 is
  -- polynomial: (0 1 2 4 5 7 8 10 11 12 16 22 23 26 32)
  -- data width: 1024
  -- convention: the first serial bit is D[1023]
  function nextCRC32_D1024
    (Data: std_logic_vector(1023 downto 0);
     crc:  std_logic_vector(31 downto 0))
    return std_logic_vector;
end PCK_CRC32_D1024;


package body PCK_CRC32_D1024 is

  -- polynomial: (0 1 2 4 5 7 8 10 11 12 16 22 23 26 32)
  -- data width: 1024
  -- convention: the first serial bit is D[1023]
  function nextCRC32_D1024
    (Data: std_logic_vector(1023 downto 0);
     crc:  std_logic_vector(31 downto 0))
    return std_logic_vector is

    variable d:      std_logic_vector(1023 downto 0);
    variable c:      std_logic_vector(31 downto 0);
    variable newcrc: std_logic_vector(31 downto 0);

  begin
    d := Data;
    c := crc;

    newcrc(0) := d(1021) xor d(1019) xor d(1018) xor d(1016) xor d(1015) xor d(1012) xor d(1011) xor d(1009) xor d(1008) xor d(1006) xor d(1005) xor d(1004) xor d(1000) xor d(999) xor d(998) xor d(996) xor d(994) xor d(992) xor d(990) xor d(985) xor d(984) xor d(983) xor d(982) xor d(981) xor d(980) xor d(979) xor d(978) xor d(977) xor d(975) xor d(974) xor d(971) xor d(967) xor d(960) xor d(959) xor d(958) xor d(955) xor d(954) xor d(953) xor d(950) xor d(948) xor d(944) xor d(941) xor d(939) xor d(938) xor d(935) xor d(934) xor d(933) xor d(931) xor d(920) xor d(918) xor d(917) xor d(915) xor d(910) xor d(907) xor d(906) xor d(904) xor d(903) xor d(902) xor d(901) xor d(900) xor d(899) xor d(898) xor d(897) xor d(896) xor d(893) xor d(891) xor d(890) xor d(889) xor d(887) xor d(886) xor d(883) xor d(881) xor d(879) xor d(878) xor d(877) xor d(876) xor d(875) xor d(874) xor d(873) xor d(871) xor d(869) xor d(868) xor d(867) xor d(863) xor d(861) xor d(860) xor d(859) xor d(857) xor d(854) xor d(853) xor d(851) xor d(850) xor d(849) xor d(848) xor d(846) xor d(842) xor d(840) xor d(839) xor d(837) xor d(835) xor d(834) xor d(832) xor d(827) xor d(825) xor d(824) xor d(819) xor d(818) xor d(816) xor d(815) xor d(814) xor d(813) xor d(812) xor d(811) xor d(810) xor d(809) xor d(808) xor d(807) xor d(806) xor d(804) xor d(803) xor d(802) xor d(800) xor d(798) xor d(793) xor d(791) xor d(788) xor d(786) xor d(785) xor d(784) xor d(782) xor d(780) xor d(776) xor d(774) xor d(769) xor d(767) xor d(765) xor d(763) xor d(762) xor d(758) xor d(756) xor d(755) xor d(753) xor d(750) xor d(748) xor d(747) xor d(744) xor d(742) xor d(741) xor d(740) xor d(736) xor d(732) xor d(731) xor d(729) xor d(727) xor d(725) xor d(724) xor d(723) xor d(722) xor d(721) xor d(720) xor d(719) xor d(715) xor d(710) xor d(708) xor d(707) xor d(704) xor d(702) xor d(701) xor d(700) xor d(698) xor d(695) xor d(694) xor d(693) xor d(691) xor d(689) xor d(687) xor d(686) xor d(680) xor d(675) xor d(674) xor d(673) xor d(672) xor d(670) xor d(669) xor d(668) xor d(667) xor d(666) xor d(665) xor d(658) xor d(656) xor d(655) xor d(653) xor d(652) xor d(649) xor d(648) xor d(646) xor d(644) xor d(642) xor d(640) xor d(636) xor d(632) xor d(630) xor d(629) xor d(626) xor d(624) xor d(623) xor d(620) xor d(619) xor d(617) xor d(615) xor d(613) xor d(612) xor d(611) xor d(610) xor d(609) xor d(607) xor d(606) xor d(604) xor d(603) xor d(602) xor d(600) xor d(599) xor d(596) xor d(595) xor d(593) xor d(592) xor d(591) xor d(587) xor d(586) xor d(585) xor d(583) xor d(580) xor d(578) xor d(575) xor d(574) xor d(573) xor d(571) xor d(567) xor d(565) xor d(563) xor d(561) xor d(560) xor d(558) xor d(557) xor d(556) xor d(555) xor d(554) xor d(551) xor d(549) xor d(545) xor d(542) xor d(540) xor d(539) xor d(535) xor d(534) xor d(532) xor d(531) xor d(530) xor d(529) xor d(528) xor d(526) xor d(525) xor d(522) xor d(521) xor d(519) xor d(518) xor d(516) xor d(514) xor d(512) xor d(511) xor d(510) xor d(508) xor d(507) xor d(506) xor d(502) xor d(501) xor d(500) xor d(495) xor d(494) xor d(493) xor d(492) xor d(491) xor d(490) xor d(489) xor d(488) xor d(486) xor d(483) xor d(482) xor d(481) xor d(480) xor d(479) xor d(477) xor d(476) xor d(472) xor d(470) xor d(468) xor d(465) xor d(464) xor d(462) xor d(461) xor d(458) xor d(452) xor d(450) xor d(449) xor d(448) xor d(444) xor d(437) xor d(436) xor d(434) xor d(433) xor d(424) xor d(422) xor d(419) xor d(418) xor d(416) xor d(414) xor d(412) xor d(409) xor d(408) xor d(407) xor d(405) xor d(404) xor d(400) xor d(399) xor d(398) xor d(396) xor d(393) xor d(392) xor d(391) xor d(390) xor d(388) xor d(387) xor d(386) xor d(381) xor d(378) xor d(376) xor d(374) xor d(372) xor d(369) xor d(368) xor d(366) xor d(363) xor d(362) xor d(359) xor d(358) xor d(357) xor d(353) xor d(349) xor d(348) xor d(347) xor d(345) xor d(344) xor d(342) xor d(341) xor d(339) xor d(338) xor d(337) xor d(335) xor d(334) xor d(333) xor d(328) xor d(327) xor d(322) xor d(321) xor d(320) xor d(319) xor d(318) xor d(317) xor d(315) xor d(312) xor d(310) xor d(309) xor d(305) xor d(303) xor d(302) xor d(300) xor d(299) xor d(298) xor d(297) xor d(296) xor d(295) xor d(294) xor d(292) xor d(290) xor d(288) xor d(287) xor d(286) xor d(283) xor d(279) xor d(277) xor d(276) xor d(274) xor d(273) xor d(269) xor d(268) xor d(265) xor d(264) xor d(261) xor d(259) xor d(257) xor d(255) xor d(252) xor d(248) xor d(243) xor d(237) xor d(234) xor d(230) xor d(228) xor d(227) xor d(226) xor d(224) xor d(216) xor d(214) xor d(212) xor d(210) xor d(209) xor d(208) xor d(207) xor d(203) xor d(202) xor d(201) xor d(199) xor d(198) xor d(197) xor d(194) xor d(193) xor d(192) xor d(191) xor d(190) xor d(188) xor d(186) xor d(183) xor d(182) xor d(172) xor d(171) xor d(170) xor d(169) xor d(167) xor d(166) xor d(162) xor d(161) xor d(158) xor d(156) xor d(155) xor d(151) xor d(149) xor d(144) xor d(143) xor d(137) xor d(136) xor d(135) xor d(134) xor d(132) xor d(128) xor d(127) xor d(126) xor d(125) xor d(123) xor d(119) xor d(118) xor d(117) xor d(116) xor d(114) xor d(113) xor d(111) xor d(110) xor d(106) xor d(104) xor d(103) xor d(101) xor d(99) xor d(98) xor d(97) xor d(96) xor d(95) xor d(94) xor d(87) xor d(85) xor d(84) xor d(83) xor d(82) xor d(81) xor d(79) xor d(73) xor d(72) xor d(68) xor d(67) xor d(66) xor d(65) xor d(63) xor d(61) xor d(60) xor d(58) xor d(55) xor d(54) xor d(53) xor d(50) xor d(48) xor d(47) xor d(45) xor d(44) xor d(37) xor d(34) xor d(32) xor d(31) xor d(30) xor d(29) xor d(28) xor d(26) xor d(25) xor d(24) xor d(16) xor d(12) xor d(10) xor d(9) xor d(6) xor d(0) xor c(0) xor c(2) xor c(4) xor c(6) xor c(7) xor c(8) xor c(12) xor c(13) xor c(14) xor c(16) xor c(17) xor c(19) xor c(20) xor c(23) xor c(24) xor c(26) xor c(27) xor c(29);
    newcrc(1) := d(1022) xor d(1021) xor d(1020) xor d(1018) xor d(1017) xor d(1015) xor d(1013) xor d(1011) xor d(1010) xor d(1008) xor d(1007) xor d(1004) xor d(1001) xor d(998) xor d(997) xor d(996) xor d(995) xor d(994) xor d(993) xor d(992) xor d(991) xor d(990) xor d(986) xor d(977) xor d(976) xor d(974) xor d(972) xor d(971) xor d(968) xor d(967) xor d(961) xor d(958) xor d(956) xor d(953) xor d(951) xor d(950) xor d(949) xor d(948) xor d(945) xor d(944) xor d(942) xor d(941) xor d(940) xor d(938) xor d(936) xor d(933) xor d(932) xor d(931) xor d(921) xor d(920) xor d(919) xor d(917) xor d(916) xor d(915) xor d(911) xor d(910) xor d(908) xor d(906) xor d(905) xor d(896) xor d(894) xor d(893) xor d(892) xor d(889) xor d(888) xor d(886) xor d(884) xor d(883) xor d(882) xor d(881) xor d(880) xor d(873) xor d(872) xor d(871) xor d(870) xor d(867) xor d(864) xor d(863) xor d(862) xor d(859) xor d(858) xor d(857) xor d(855) xor d(853) xor d(852) xor d(848) xor d(847) xor d(846) xor d(843) xor d(842) xor d(841) xor d(839) xor d(838) xor d(837) xor d(836) xor d(834) xor d(833) xor d(832) xor d(828) xor d(827) xor d(826) xor d(824) xor d(820) xor d(818) xor d(817) xor d(806) xor d(805) xor d(802) xor d(801) xor d(800) xor d(799) xor d(798) xor d(794) xor d(793) xor d(792) xor d(791) xor d(789) xor d(788) xor d(787) xor d(784) xor d(783) xor d(782) xor d(781) xor d(780) xor d(777) xor d(776) xor d(775) xor d(774) xor d(770) xor d(769) xor d(768) xor d(767) xor d(766) xor d(765) xor d(764) xor d(762) xor d(759) xor d(758) xor d(757) xor d(755) xor d(754) xor d(753) xor d(751) xor d(750) xor d(749) xor d(747) xor d(745) xor d(744) xor d(743) xor d(740) xor d(737) xor d(736) xor d(733) xor d(731) xor d(730) xor d(729) xor d(728) xor d(727) xor d(726) xor d(719) xor d(716) xor d(715) xor d(711) xor d(710) xor d(709) xor d(707) xor d(705) xor d(704) xor d(703) xor d(700) xor d(699) xor d(698) xor d(696) xor d(693) xor d(692) xor d(691) xor d(690) xor d(689) xor d(688) xor d(686) xor d(681) xor d(680) xor d(676) xor d(672) xor d(671) xor d(665) xor d(659) xor d(658) xor d(657) xor d(655) xor d(654) xor d(652) xor d(650) xor d(648) xor d(647) xor d(646) xor d(645) xor d(644) xor d(643) xor d(642) xor d(641) xor d(640) xor d(637) xor d(636) xor d(633) xor d(632) xor d(631) xor d(629) xor d(627) xor d(626) xor d(625) xor d(623) xor d(621) xor d(619) xor d(618) xor d(617) xor d(616) xor d(615) xor d(614) xor d(609) xor d(608) xor d(606) xor d(605) xor d(602) xor d(601) xor d(599) xor d(597) xor d(595) xor d(594) xor d(591) xor d(588) xor d(585) xor d(584) xor d(583) xor d(581) xor d(580) xor d(579) xor d(578) xor d(576) xor d(573) xor d(572) xor d(571) xor d(568) xor d(567) xor d(566) xor d(565) xor d(564) xor d(563) xor d(562) xor d(560) xor d(559) xor d(554) xor d(552) xor d(551) xor d(550) xor d(549) xor d(546) xor d(545) xor d(543) xor d(542) xor d(541) xor d(539) xor d(536) xor d(534) xor d(533) xor d(528) xor d(527) xor d(525) xor d(523) xor d(521) xor d(520) xor d(518) xor d(517) xor d(516) xor d(515) xor d(514) xor d(513) xor d(510) xor d(509) xor d(506) xor d(503) xor d(500) xor d(496) xor d(488) xor d(487) xor d(486) xor d(484) xor d(479) xor d(478) xor d(476) xor d(473) xor d(472) xor d(471) xor d(470) xor d(469) xor d(468) xor d(466) xor d(464) xor d(463) xor d(461) xor d(459) xor d(458) xor d(453) xor d(452) xor d(451) xor d(448) xor d(445) xor d(444) xor d(438) xor d(436) xor d(435) xor d(433) xor d(425) xor d(424) xor d(423) xor d(422) xor d(420) xor d(418) xor d(417) xor d(416) xor d(415) xor d(414) xor d(413) xor d(412) xor d(410) xor d(407) xor d(406) xor d(404) xor d(401) xor d(398) xor d(397) xor d(396) xor d(394) xor d(390) xor d(389) xor d(386) xor d(382) xor d(381) xor d(379) xor d(378) xor d(377) xor d(376) xor d(375) xor d(374) xor d(373) xor d(372) xor d(370) xor d(368) xor d(367) xor d(366) xor d(364) xor d(362) xor d(360) xor d(357) xor d(354) xor d(353) xor d(350) xor d(347) xor d(346) xor d(344) xor d(343) xor d(341) xor d(340) xor d(337) xor d(336) xor d(333) xor d(329) xor d(327) xor d(323) xor d(317) xor d(316) xor d(315) xor d(313) xor d(312) xor d(311) xor d(309) xor d(306) xor d(305) xor d(304) xor d(302) xor d(301) xor d(294) xor d(293) xor d(292) xor d(291) xor d(290) xor d(289) xor d(286) xor d(284) xor d(283) xor d(280) xor d(279) xor d(278) xor d(276) xor d(275) xor d(273) xor d(270) xor d(268) xor d(266) xor d(264) xor d(262) xor d(261) xor d(260) xor d(259) xor d(258) xor d(257) xor d(256) xor d(255) xor d(253) xor d(252) xor d(249) xor d(248) xor d(244) xor d(243) xor d(238) xor d(237) xor d(235) xor d(234) xor d(231) xor d(230) xor d(229) xor d(226) xor d(225) xor d(224) xor d(217) xor d(216) xor d(215) xor d(214) xor d(213) xor d(212) xor d(211) xor d(207) xor d(204) xor d(201) xor d(200) xor d(197) xor d(195) xor d(190) xor d(189) xor d(188) xor d(187) xor d(186) xor d(184) xor d(182) xor d(173) xor d(169) xor d(168) xor d(166) xor d(163) xor d(161) xor d(159) xor d(158) xor d(157) xor d(155) xor d(152) xor d(151) xor d(150) xor d(149) xor d(145) xor d(143) xor d(138) xor d(134) xor d(133) xor d(132) xor d(129) xor d(125) xor d(124) xor d(123) xor d(120) xor d(116) xor d(115) xor d(113) xor d(112) xor d(110) xor d(107) xor d(106) xor d(105) xor d(103) xor d(102) xor d(101) xor d(100) xor d(94) xor d(88) xor d(87) xor d(86) xor d(81) xor d(80) xor d(79) xor d(74) xor d(72) xor d(69) xor d(65) xor d(64) xor d(63) xor d(62) xor d(60) xor d(59) xor d(58) xor d(56) xor d(53) xor d(51) xor d(50) xor d(49) xor d(47) xor d(46) xor d(44) xor d(38) xor d(37) xor d(35) xor d(34) xor d(33) xor d(28) xor d(27) xor d(24) xor d(17) xor d(16) xor d(13) xor d(12) xor d(11) xor d(9) xor d(7) xor d(6) xor d(1) xor d(0) xor c(0) xor c(1) xor c(2) xor c(3) xor c(4) xor c(5) xor c(6) xor c(9) xor c(12) xor c(15) xor c(16) xor c(18) xor c(19) xor c(21) xor c(23) xor c(25) xor c(26) xor c(28) xor c(29) xor c(30);
    newcrc(2) := d(1023) xor d(1022) xor d(1015) xor d(1014) xor d(1006) xor d(1004) xor d(1002) xor d(1000) xor d(997) xor d(995) xor d(993) xor d(991) xor d(990) xor d(987) xor d(985) xor d(984) xor d(983) xor d(982) xor d(981) xor d(980) xor d(979) xor d(974) xor d(973) xor d(972) xor d(971) xor d(969) xor d(968) xor d(967) xor d(962) xor d(960) xor d(958) xor d(957) xor d(955) xor d(953) xor d(952) xor d(951) xor d(949) xor d(948) xor d(946) xor d(945) xor d(944) xor d(943) xor d(942) xor d(938) xor d(937) xor d(935) xor d(932) xor d(931) xor d(922) xor d(921) xor d(916) xor d(915) xor d(912) xor d(911) xor d(910) xor d(909) xor d(904) xor d(903) xor d(902) xor d(901) xor d(900) xor d(899) xor d(898) xor d(896) xor d(895) xor d(894) xor d(891) xor d(886) xor d(885) xor d(884) xor d(882) xor d(879) xor d(878) xor d(877) xor d(876) xor d(875) xor d(872) xor d(869) xor d(867) xor d(865) xor d(864) xor d(861) xor d(858) xor d(857) xor d(856) xor d(851) xor d(850) xor d(847) xor d(846) xor d(844) xor d(843) xor d(838) xor d(833) xor d(832) xor d(829) xor d(828) xor d(824) xor d(821) xor d(816) xor d(815) xor d(814) xor d(813) xor d(812) xor d(811) xor d(810) xor d(809) xor d(808) xor d(804) xor d(801) xor d(799) xor d(798) xor d(795) xor d(794) xor d(792) xor d(791) xor d(790) xor d(789) xor d(786) xor d(783) xor d(781) xor d(780) xor d(778) xor d(777) xor d(775) xor d(774) xor d(771) xor d(770) xor d(768) xor d(766) xor d(762) xor d(760) xor d(759) xor d(754) xor d(753) xor d(752) xor d(751) xor d(747) xor d(746) xor d(745) xor d(742) xor d(740) xor d(738) xor d(737) xor d(736) xor d(734) xor d(730) xor d(728) xor d(725) xor d(724) xor d(723) xor d(722) xor d(721) xor d(719) xor d(717) xor d(716) xor d(715) xor d(712) xor d(711) xor d(707) xor d(706) xor d(705) xor d(702) xor d(699) xor d(698) xor d(697) xor d(695) xor d(692) xor d(690) xor d(686) xor d(682) xor d(681) xor d(680) xor d(677) xor d(675) xor d(674) xor d(670) xor d(669) xor d(668) xor d(667) xor d(665) xor d(660) xor d(659) xor d(652) xor d(651) xor d(647) xor d(645) xor d(643) xor d(641) xor d(640) xor d(638) xor d(637) xor d(636) xor d(634) xor d(633) xor d(629) xor d(628) xor d(627) xor d(623) xor d(622) xor d(618) xor d(616) xor d(613) xor d(612) xor d(611) xor d(604) xor d(599) xor d(598) xor d(593) xor d(591) xor d(589) xor d(587) xor d(584) xor d(583) xor d(582) xor d(581) xor d(579) xor d(578) xor d(577) xor d(575) xor d(572) xor d(571) xor d(569) xor d(568) xor d(566) xor d(564) xor d(558) xor d(557) xor d(556) xor d(554) xor d(553) xor d(552) xor d(550) xor d(549) xor d(547) xor d(546) xor d(545) xor d(544) xor d(543) xor d(539) xor d(537) xor d(532) xor d(531) xor d(530) xor d(525) xor d(524) xor d(517) xor d(515) xor d(512) xor d(508) xor d(506) xor d(504) xor d(502) xor d(500) xor d(497) xor d(495) xor d(494) xor d(493) xor d(492) xor d(491) xor d(490) xor d(487) xor d(486) xor d(485) xor d(483) xor d(482) xor d(481) xor d(476) xor d(474) xor d(473) xor d(471) xor d(469) xor d(468) xor d(467) xor d(461) xor d(460) xor d(459) xor d(458) xor d(454) xor d(453) xor d(450) xor d(448) xor d(446) xor d(445) xor d(444) xor d(439) xor d(433) xor d(426) xor d(425) xor d(423) xor d(422) xor d(421) xor d(417) xor d(415) xor d(413) xor d(412) xor d(411) xor d(409) xor d(404) xor d(402) xor d(400) xor d(397) xor d(396) xor d(395) xor d(393) xor d(392) xor d(388) xor d(386) xor d(383) xor d(382) xor d(381) xor d(380) xor d(379) xor d(377) xor d(375) xor d(373) xor d(372) xor d(371) xor d(367) xor d(366) xor d(365) xor d(362) xor d(361) xor d(359) xor d(357) xor d(355) xor d(354) xor d(353) xor d(351) xor d(349) xor d(339) xor d(335) xor d(333) xor d(330) xor d(327) xor d(324) xor d(322) xor d(321) xor d(320) xor d(319) xor d(316) xor d(315) xor d(314) xor d(313) xor d(309) xor d(307) xor d(306) xor d(300) xor d(299) xor d(298) xor d(297) xor d(296) xor d(293) xor d(291) xor d(288) xor d(286) xor d(285) xor d(284) xor d(283) xor d(281) xor d(280) xor d(273) xor d(271) xor d(268) xor d(267) xor d(264) xor d(263) xor d(262) xor d(260) xor d(258) xor d(256) xor d(255) xor d(254) xor d(253) xor d(252) xor d(250) xor d(249) xor d(248) xor d(245) xor d(244) xor d(243) xor d(239) xor d(238) xor d(237) xor d(236) xor d(235) xor d(234) xor d(232) xor d(231) xor d(228) xor d(225) xor d(224) xor d(218) xor d(217) xor d(215) xor d(213) xor d(210) xor d(209) xor d(207) xor d(205) xor d(203) xor d(199) xor d(197) xor d(196) xor d(194) xor d(193) xor d(192) xor d(189) xor d(187) xor d(186) xor d(185) xor d(182) xor d(174) xor d(172) xor d(171) xor d(166) xor d(164) xor d(161) xor d(160) xor d(159) xor d(155) xor d(153) xor d(152) xor d(150) xor d(149) xor d(146) xor d(143) xor d(139) xor d(137) xor d(136) xor d(133) xor d(132) xor d(130) xor d(128) xor d(127) xor d(124) xor d(123) xor d(121) xor d(119) xor d(118) xor d(110) xor d(108) xor d(107) xor d(102) xor d(99) xor d(98) xor d(97) xor d(96) xor d(94) xor d(89) xor d(88) xor d(85) xor d(84) xor d(83) xor d(80) xor d(79) xor d(75) xor d(72) xor d(70) xor d(68) xor d(67) xor d(64) xor d(59) xor d(58) xor d(57) xor d(55) xor d(53) xor d(52) xor d(51) xor d(44) xor d(39) xor d(38) xor d(37) xor d(36) xor d(35) xor d(32) xor d(31) xor d(30) xor d(26) xor d(24) xor d(18) xor d(17) xor d(16) xor d(14) xor d(13) xor d(9) xor d(8) xor d(7) xor d(6) xor d(2) xor d(1) xor d(0) xor c(1) xor c(3) xor c(5) xor c(8) xor c(10) xor c(12) xor c(14) xor c(22) xor c(23) xor c(30) xor c(31);
    newcrc(3) := d(1023) xor d(1016) xor d(1015) xor d(1007) xor d(1005) xor d(1003) xor d(1001) xor d(998) xor d(996) xor d(994) xor d(992) xor d(991) xor d(988) xor d(986) xor d(985) xor d(984) xor d(983) xor d(982) xor d(981) xor d(980) xor d(975) xor d(974) xor d(973) xor d(972) xor d(970) xor d(969) xor d(968) xor d(963) xor d(961) xor d(959) xor d(958) xor d(956) xor d(954) xor d(953) xor d(952) xor d(950) xor d(949) xor d(947) xor d(946) xor d(945) xor d(944) xor d(943) xor d(939) xor d(938) xor d(936) xor d(933) xor d(932) xor d(923) xor d(922) xor d(917) xor d(916) xor d(913) xor d(912) xor d(911) xor d(910) xor d(905) xor d(904) xor d(903) xor d(902) xor d(901) xor d(900) xor d(899) xor d(897) xor d(896) xor d(895) xor d(892) xor d(887) xor d(886) xor d(885) xor d(883) xor d(880) xor d(879) xor d(878) xor d(877) xor d(876) xor d(873) xor d(870) xor d(868) xor d(866) xor d(865) xor d(862) xor d(859) xor d(858) xor d(857) xor d(852) xor d(851) xor d(848) xor d(847) xor d(845) xor d(844) xor d(839) xor d(834) xor d(833) xor d(830) xor d(829) xor d(825) xor d(822) xor d(817) xor d(816) xor d(815) xor d(814) xor d(813) xor d(812) xor d(811) xor d(810) xor d(809) xor d(805) xor d(802) xor d(800) xor d(799) xor d(796) xor d(795) xor d(793) xor d(792) xor d(791) xor d(790) xor d(787) xor d(784) xor d(782) xor d(781) xor d(779) xor d(778) xor d(776) xor d(775) xor d(772) xor d(771) xor d(769) xor d(767) xor d(763) xor d(761) xor d(760) xor d(755) xor d(754) xor d(753) xor d(752) xor d(748) xor d(747) xor d(746) xor d(743) xor d(741) xor d(739) xor d(738) xor d(737) xor d(735) xor d(731) xor d(729) xor d(726) xor d(725) xor d(724) xor d(723) xor d(722) xor d(720) xor d(718) xor d(717) xor d(716) xor d(713) xor d(712) xor d(708) xor d(707) xor d(706) xor d(703) xor d(700) xor d(699) xor d(698) xor d(696) xor d(693) xor d(691) xor d(687) xor d(683) xor d(682) xor d(681) xor d(678) xor d(676) xor d(675) xor d(671) xor d(670) xor d(669) xor d(668) xor d(666) xor d(661) xor d(660) xor d(653) xor d(652) xor d(648) xor d(646) xor d(644) xor d(642) xor d(641) xor d(639) xor d(638) xor d(637) xor d(635) xor d(634) xor d(630) xor d(629) xor d(628) xor d(624) xor d(623) xor d(619) xor d(617) xor d(614) xor d(613) xor d(612) xor d(605) xor d(600) xor d(599) xor d(594) xor d(592) xor d(590) xor d(588) xor d(585) xor d(584) xor d(583) xor d(582) xor d(580) xor d(579) xor d(578) xor d(576) xor d(573) xor d(572) xor d(570) xor d(569) xor d(567) xor d(565) xor d(559) xor d(558) xor d(557) xor d(555) xor d(554) xor d(553) xor d(551) xor d(550) xor d(548) xor d(547) xor d(546) xor d(545) xor d(544) xor d(540) xor d(538) xor d(533) xor d(532) xor d(531) xor d(526) xor d(525) xor d(518) xor d(516) xor d(513) xor d(509) xor d(507) xor d(505) xor d(503) xor d(501) xor d(498) xor d(496) xor d(495) xor d(494) xor d(493) xor d(492) xor d(491) xor d(488) xor d(487) xor d(486) xor d(484) xor d(483) xor d(482) xor d(477) xor d(475) xor d(474) xor d(472) xor d(470) xor d(469) xor d(468) xor d(462) xor d(461) xor d(460) xor d(459) xor d(455) xor d(454) xor d(451) xor d(449) xor d(447) xor d(446) xor d(445) xor d(440) xor d(434) xor d(427) xor d(426) xor d(424) xor d(423) xor d(422) xor d(418) xor d(416) xor d(414) xor d(413) xor d(412) xor d(410) xor d(405) xor d(403) xor d(401) xor d(398) xor d(397) xor d(396) xor d(394) xor d(393) xor d(389) xor d(387) xor d(384) xor d(383) xor d(382) xor d(381) xor d(380) xor d(378) xor d(376) xor d(374) xor d(373) xor d(372) xor d(368) xor d(367) xor d(366) xor d(363) xor d(362) xor d(360) xor d(358) xor d(356) xor d(355) xor d(354) xor d(352) xor d(350) xor d(340) xor d(336) xor d(334) xor d(331) xor d(328) xor d(325) xor d(323) xor d(322) xor d(321) xor d(320) xor d(317) xor d(316) xor d(315) xor d(314) xor d(310) xor d(308) xor d(307) xor d(301) xor d(300) xor d(299) xor d(298) xor d(297) xor d(294) xor d(292) xor d(289) xor d(287) xor d(286) xor d(285) xor d(284) xor d(282) xor d(281) xor d(274) xor d(272) xor d(269) xor d(268) xor d(265) xor d(264) xor d(263) xor d(261) xor d(259) xor d(257) xor d(256) xor d(255) xor d(254) xor d(253) xor d(251) xor d(250) xor d(249) xor d(246) xor d(245) xor d(244) xor d(240) xor d(239) xor d(238) xor d(237) xor d(236) xor d(235) xor d(233) xor d(232) xor d(229) xor d(226) xor d(225) xor d(219) xor d(218) xor d(216) xor d(214) xor d(211) xor d(210) xor d(208) xor d(206) xor d(204) xor d(200) xor d(198) xor d(197) xor d(195) xor d(194) xor d(193) xor d(190) xor d(188) xor d(187) xor d(186) xor d(183) xor d(175) xor d(173) xor d(172) xor d(167) xor d(165) xor d(162) xor d(161) xor d(160) xor d(156) xor d(154) xor d(153) xor d(151) xor d(150) xor d(147) xor d(144) xor d(140) xor d(138) xor d(137) xor d(134) xor d(133) xor d(131) xor d(129) xor d(128) xor d(125) xor d(124) xor d(122) xor d(120) xor d(119) xor d(111) xor d(109) xor d(108) xor d(103) xor d(100) xor d(99) xor d(98) xor d(97) xor d(95) xor d(90) xor d(89) xor d(86) xor d(85) xor d(84) xor d(81) xor d(80) xor d(76) xor d(73) xor d(71) xor d(69) xor d(68) xor d(65) xor d(60) xor d(59) xor d(58) xor d(56) xor d(54) xor d(53) xor d(52) xor d(45) xor d(40) xor d(39) xor d(38) xor d(37) xor d(36) xor d(33) xor d(32) xor d(31) xor d(27) xor d(25) xor d(19) xor d(18) xor d(17) xor d(15) xor d(14) xor d(10) xor d(9) xor d(8) xor d(7) xor d(3) xor d(2) xor d(1) xor c(0) xor c(2) xor c(4) xor c(6) xor c(9) xor c(11) xor c(13) xor c(15) xor c(23) xor c(24) xor c(31);
    newcrc(4) := d(1021) xor d(1019) xor d(1018) xor d(1017) xor d(1015) xor d(1012) xor d(1011) xor d(1009) xor d(1005) xor d(1002) xor d(1000) xor d(998) xor d(997) xor d(996) xor d(995) xor d(994) xor d(993) xor d(990) xor d(989) xor d(987) xor d(986) xor d(980) xor d(979) xor d(978) xor d(977) xor d(976) xor d(973) xor d(970) xor d(969) xor d(967) xor d(964) xor d(962) xor d(958) xor d(957) xor d(951) xor d(947) xor d(946) xor d(945) xor d(941) xor d(940) xor d(938) xor d(937) xor d(935) xor d(931) xor d(924) xor d(923) xor d(920) xor d(915) xor d(914) xor d(913) xor d(912) xor d(911) xor d(910) xor d(907) xor d(905) xor d(899) xor d(891) xor d(890) xor d(889) xor d(888) xor d(884) xor d(883) xor d(880) xor d(876) xor d(875) xor d(873) xor d(868) xor d(866) xor d(861) xor d(858) xor d(857) xor d(854) xor d(852) xor d(851) xor d(850) xor d(845) xor d(842) xor d(839) xor d(837) xor d(832) xor d(831) xor d(830) xor d(827) xor d(826) xor d(825) xor d(824) xor d(823) xor d(819) xor d(817) xor d(809) xor d(808) xor d(807) xor d(804) xor d(802) xor d(801) xor d(798) xor d(797) xor d(796) xor d(794) xor d(792) xor d(786) xor d(784) xor d(783) xor d(779) xor d(777) xor d(774) xor d(773) xor d(772) xor d(770) xor d(769) xor d(768) xor d(767) xor d(765) xor d(764) xor d(763) xor d(761) xor d(758) xor d(754) xor d(750) xor d(749) xor d(741) xor d(739) xor d(738) xor d(731) xor d(730) xor d(729) xor d(726) xor d(722) xor d(720) xor d(718) xor d(717) xor d(715) xor d(714) xor d(713) xor d(710) xor d(709) xor d(702) xor d(699) xor d(698) xor d(697) xor d(695) xor d(693) xor d(692) xor d(691) xor d(689) xor d(688) xor d(687) xor d(686) xor d(684) xor d(683) xor d(682) xor d(680) xor d(679) xor d(677) xor d(676) xor d(675) xor d(674) xor d(673) xor d(671) xor d(668) xor d(666) xor d(665) xor d(662) xor d(661) xor d(658) xor d(656) xor d(655) xor d(654) xor d(652) xor d(648) xor d(647) xor d(646) xor d(645) xor d(644) xor d(643) xor d(639) xor d(638) xor d(635) xor d(632) xor d(631) xor d(626) xor d(625) xor d(623) xor d(619) xor d(618) xor d(617) xor d(614) xor d(612) xor d(611) xor d(610) xor d(609) xor d(607) xor d(604) xor d(603) xor d(602) xor d(601) xor d(599) xor d(596) xor d(592) xor d(589) xor d(587) xor d(584) xor d(581) xor d(579) xor d(578) xor d(577) xor d(575) xor d(570) xor d(568) xor d(567) xor d(566) xor d(565) xor d(563) xor d(561) xor d(559) xor d(557) xor d(552) xor d(548) xor d(547) xor d(546) xor d(542) xor d(541) xor d(540) xor d(535) xor d(533) xor d(531) xor d(530) xor d(529) xor d(528) xor d(527) xor d(525) xor d(522) xor d(521) xor d(518) xor d(517) xor d(516) xor d(512) xor d(511) xor d(507) xor d(504) xor d(501) xor d(500) xor d(499) xor d(497) xor d(496) xor d(491) xor d(490) xor d(487) xor d(486) xor d(485) xor d(484) xor d(482) xor d(481) xor d(480) xor d(479) xor d(478) xor d(477) xor d(475) xor d(473) xor d(472) xor d(471) xor d(469) xor d(468) xor d(465) xor d(464) xor d(463) xor d(460) xor d(458) xor d(456) xor d(455) xor d(449) xor d(447) xor d(446) xor d(444) xor d(441) xor d(437) xor d(436) xor d(435) xor d(434) xor d(433) xor d(428) xor d(427) xor d(425) xor d(423) xor d(422) xor d(418) xor d(417) xor d(416) xor d(415) xor d(413) xor d(412) xor d(411) xor d(409) xor d(408) xor d(407) xor d(406) xor d(405) xor d(402) xor d(400) xor d(397) xor d(396) xor d(395) xor d(394) xor d(393) xor d(392) xor d(391) xor d(387) xor d(386) xor d(385) xor d(384) xor d(383) xor d(382) xor d(379) xor d(378) xor d(377) xor d(376) xor d(375) xor d(373) xor d(372) xor d(367) xor d(366) xor d(364) xor d(362) xor d(361) xor d(358) xor d(356) xor d(355) xor d(351) xor d(349) xor d(348) xor d(347) xor d(345) xor d(344) xor d(342) xor d(339) xor d(338) xor d(334) xor d(333) xor d(332) xor d(329) xor d(328) xor d(327) xor d(326) xor d(324) xor d(323) xor d(320) xor d(319) xor d(316) xor d(312) xor d(311) xor d(310) xor d(308) xor d(305) xor d(303) xor d(301) xor d(297) xor d(296) xor d(294) xor d(293) xor d(292) xor d(285) xor d(282) xor d(279) xor d(277) xor d(276) xor d(275) xor d(274) xor d(270) xor d(268) xor d(266) xor d(262) xor d(261) xor d(260) xor d(259) xor d(258) xor d(256) xor d(254) xor d(251) xor d(250) xor d(248) xor d(247) xor d(246) xor d(245) xor d(243) xor d(241) xor d(240) xor d(239) xor d(238) xor d(236) xor d(233) xor d(228) xor d(224) xor d(220) xor d(219) xor d(217) xor d(216) xor d(215) xor d(214) xor d(211) xor d(210) xor d(208) xor d(205) xor d(203) xor d(202) xor d(197) xor d(196) xor d(195) xor d(193) xor d(192) xor d(190) xor d(189) xor d(187) xor d(186) xor d(184) xor d(183) xor d(182) xor d(176) xor d(174) xor d(173) xor d(172) xor d(171) xor d(170) xor d(169) xor d(168) xor d(167) xor d(163) xor d(158) xor d(157) xor d(156) xor d(154) xor d(152) xor d(149) xor d(148) xor d(145) xor d(144) xor d(143) xor d(141) xor d(139) xor d(138) xor d(137) xor d(136) xor d(130) xor d(129) xor d(128) xor d(127) xor d(121) xor d(120) xor d(119) xor d(118) xor d(117) xor d(116) xor d(114) xor d(113) xor d(112) xor d(111) xor d(109) xor d(106) xor d(103) xor d(100) xor d(97) xor d(95) xor d(94) xor d(91) xor d(90) xor d(86) xor d(84) xor d(83) xor d(79) xor d(77) xor d(74) xor d(73) xor d(70) xor d(69) xor d(68) xor d(67) xor d(65) xor d(63) xor d(59) xor d(58) xor d(57) xor d(50) xor d(48) xor d(47) xor d(46) xor d(45) xor d(44) xor d(41) xor d(40) xor d(39) xor d(38) xor d(33) xor d(31) xor d(30) xor d(29) xor d(25) xor d(24) xor d(20) xor d(19) xor d(18) xor d(15) xor d(12) xor d(11) xor d(8) xor d(6) xor d(4) xor d(3) xor d(2) xor d(0) xor c(1) xor c(2) xor c(3) xor c(4) xor c(5) xor c(6) xor c(8) xor c(10) xor c(13) xor c(17) xor c(19) xor c(20) xor c(23) xor c(25) xor c(26) xor c(27) xor c(29);
    newcrc(5) := d(1022) xor d(1021) xor d(1020) xor d(1015) xor d(1013) xor d(1011) xor d(1010) xor d(1009) xor d(1008) xor d(1005) xor d(1004) xor d(1003) xor d(1001) xor d(1000) xor d(997) xor d(995) xor d(992) xor d(991) xor d(988) xor d(987) xor d(985) xor d(984) xor d(983) xor d(982) xor d(975) xor d(970) xor d(968) xor d(967) xor d(965) xor d(963) xor d(960) xor d(955) xor d(954) xor d(953) xor d(952) xor d(950) xor d(947) xor d(946) xor d(944) xor d(942) xor d(936) xor d(935) xor d(934) xor d(933) xor d(932) xor d(931) xor d(925) xor d(924) xor d(921) xor d(920) xor d(918) xor d(917) xor d(916) xor d(914) xor d(913) xor d(912) xor d(911) xor d(910) xor d(908) xor d(907) xor d(904) xor d(903) xor d(902) xor d(901) xor d(899) xor d(898) xor d(897) xor d(896) xor d(893) xor d(892) xor d(887) xor d(886) xor d(885) xor d(884) xor d(883) xor d(879) xor d(878) xor d(875) xor d(873) xor d(871) xor d(868) xor d(863) xor d(862) xor d(861) xor d(860) xor d(858) xor d(857) xor d(855) xor d(854) xor d(852) xor d(850) xor d(849) xor d(848) xor d(843) xor d(842) xor d(839) xor d(838) xor d(837) xor d(835) xor d(834) xor d(833) xor d(831) xor d(828) xor d(826) xor d(820) xor d(819) xor d(816) xor d(815) xor d(814) xor d(813) xor d(812) xor d(811) xor d(807) xor d(806) xor d(805) xor d(804) xor d(800) xor d(799) xor d(797) xor d(795) xor d(791) xor d(788) xor d(787) xor d(786) xor d(782) xor d(778) xor d(776) xor d(775) xor d(773) xor d(771) xor d(770) xor d(768) xor d(767) xor d(766) xor d(764) xor d(763) xor d(759) xor d(758) xor d(756) xor d(753) xor d(751) xor d(748) xor d(747) xor d(744) xor d(741) xor d(739) xor d(736) xor d(730) xor d(729) xor d(725) xor d(724) xor d(722) xor d(720) xor d(718) xor d(716) xor d(714) xor d(711) xor d(708) xor d(707) xor d(704) xor d(703) xor d(702) xor d(701) xor d(699) xor d(696) xor d(695) xor d(692) xor d(691) xor d(690) xor d(688) xor d(686) xor d(685) xor d(684) xor d(683) xor d(681) xor d(678) xor d(677) xor d(676) xor d(673) xor d(670) xor d(668) xor d(665) xor d(663) xor d(662) xor d(659) xor d(658) xor d(657) xor d(652) xor d(647) xor d(645) xor d(642) xor d(639) xor d(633) xor d(630) xor d(629) xor d(627) xor d(623) xor d(618) xor d(617) xor d(609) xor d(608) xor d(607) xor d(606) xor d(605) xor d(599) xor d(597) xor d(596) xor d(595) xor d(592) xor d(591) xor d(590) xor d(588) xor d(587) xor d(586) xor d(583) xor d(582) xor d(579) xor d(576) xor d(575) xor d(574) xor d(573) xor d(569) xor d(568) xor d(566) xor d(565) xor d(564) xor d(563) xor d(562) xor d(561) xor d(557) xor d(556) xor d(555) xor d(554) xor d(553) xor d(551) xor d(548) xor d(547) xor d(545) xor d(543) xor d(541) xor d(540) xor d(539) xor d(536) xor d(535) xor d(525) xor d(523) xor d(521) xor d(517) xor d(516) xor d(514) xor d(513) xor d(511) xor d(510) xor d(507) xor d(506) xor d(505) xor d(498) xor d(497) xor d(495) xor d(494) xor d(493) xor d(490) xor d(489) xor d(487) xor d(485) xor d(478) xor d(477) xor d(474) xor d(473) xor d(469) xor d(468) xor d(466) xor d(462) xor d(459) xor d(458) xor d(457) xor d(456) xor d(452) xor d(449) xor d(447) xor d(445) xor d(444) xor d(442) xor d(438) xor d(435) xor d(433) xor d(429) xor d(428) xor d(426) xor d(423) xor d(422) xor d(417) xor d(413) xor d(410) xor d(406) xor d(405) xor d(404) xor d(403) xor d(401) xor d(400) xor d(399) xor d(397) xor d(395) xor d(394) xor d(391) xor d(390) xor d(385) xor d(384) xor d(383) xor d(381) xor d(380) xor d(379) xor d(377) xor d(373) xor d(372) xor d(369) xor d(367) xor d(366) xor d(365) xor d(358) xor d(356) xor d(353) xor d(352) xor d(350) xor d(347) xor d(346) xor d(344) xor d(343) xor d(342) xor d(341) xor d(340) xor d(338) xor d(337) xor d(330) xor d(329) xor d(325) xor d(324) xor d(322) xor d(319) xor d(318) xor d(315) xor d(313) xor d(311) xor d(310) xor d(306) xor d(305) xor d(304) xor d(303) xor d(300) xor d(299) xor d(296) xor d(293) xor d(292) xor d(290) xor d(288) xor d(287) xor d(280) xor d(279) xor d(278) xor d(275) xor d(274) xor d(273) xor d(271) xor d(268) xor d(267) xor d(265) xor d(264) xor d(263) xor d(262) xor d(260) xor d(251) xor d(249) xor d(247) xor d(246) xor d(244) xor d(243) xor d(242) xor d(241) xor d(240) xor d(239) xor d(230) xor d(229) xor d(228) xor d(227) xor d(226) xor d(225) xor d(224) xor d(221) xor d(220) xor d(218) xor d(217) xor d(215) xor d(214) xor d(211) xor d(210) xor d(208) xor d(207) xor d(206) xor d(204) xor d(202) xor d(201) xor d(199) xor d(196) xor d(192) xor d(187) xor d(186) xor d(185) xor d(184) xor d(182) xor d(177) xor d(175) xor d(174) xor d(173) xor d(168) xor d(167) xor d(166) xor d(164) xor d(162) xor d(161) xor d(159) xor d(157) xor d(156) xor d(153) xor d(151) xor d(150) xor d(146) xor d(145) xor d(143) xor d(142) xor d(140) xor d(139) xor d(138) xor d(136) xor d(135) xor d(134) xor d(132) xor d(131) xor d(130) xor d(129) xor d(127) xor d(126) xor d(125) xor d(123) xor d(122) xor d(121) xor d(120) xor d(116) xor d(115) xor d(112) xor d(111) xor d(107) xor d(106) xor d(103) xor d(99) xor d(97) xor d(94) xor d(92) xor d(91) xor d(83) xor d(82) xor d(81) xor d(80) xor d(79) xor d(78) xor d(75) xor d(74) xor d(73) xor d(72) xor d(71) xor d(70) xor d(69) xor d(67) xor d(65) xor d(64) xor d(63) xor d(61) xor d(59) xor d(55) xor d(54) xor d(53) xor d(51) xor d(50) xor d(49) xor d(46) xor d(44) xor d(42) xor d(41) xor d(40) xor d(39) xor d(37) xor d(29) xor d(28) xor d(24) xor d(21) xor d(20) xor d(19) xor d(13) xor d(10) xor d(7) xor d(6) xor d(5) xor d(4) xor d(3) xor d(1) xor d(0) xor c(0) xor c(3) xor c(5) xor c(8) xor c(9) xor c(11) xor c(12) xor c(13) xor c(16) xor c(17) xor c(18) xor c(19) xor c(21) xor c(23) xor c(28) xor c(29) xor c(30);
    newcrc(6) := d(1023) xor d(1022) xor d(1021) xor d(1016) xor d(1014) xor d(1012) xor d(1011) xor d(1010) xor d(1009) xor d(1006) xor d(1005) xor d(1004) xor d(1002) xor d(1001) xor d(998) xor d(996) xor d(993) xor d(992) xor d(989) xor d(988) xor d(986) xor d(985) xor d(984) xor d(983) xor d(976) xor d(971) xor d(969) xor d(968) xor d(966) xor d(964) xor d(961) xor d(956) xor d(955) xor d(954) xor d(953) xor d(951) xor d(948) xor d(947) xor d(945) xor d(943) xor d(937) xor d(936) xor d(935) xor d(934) xor d(933) xor d(932) xor d(926) xor d(925) xor d(922) xor d(921) xor d(919) xor d(918) xor d(917) xor d(915) xor d(914) xor d(913) xor d(912) xor d(911) xor d(909) xor d(908) xor d(905) xor d(904) xor d(903) xor d(902) xor d(900) xor d(899) xor d(898) xor d(897) xor d(894) xor d(893) xor d(888) xor d(887) xor d(886) xor d(885) xor d(884) xor d(880) xor d(879) xor d(876) xor d(874) xor d(872) xor d(869) xor d(864) xor d(863) xor d(862) xor d(861) xor d(859) xor d(858) xor d(856) xor d(855) xor d(853) xor d(851) xor d(850) xor d(849) xor d(844) xor d(843) xor d(840) xor d(839) xor d(838) xor d(836) xor d(835) xor d(834) xor d(832) xor d(829) xor d(827) xor d(821) xor d(820) xor d(817) xor d(816) xor d(815) xor d(814) xor d(813) xor d(812) xor d(808) xor d(807) xor d(806) xor d(805) xor d(801) xor d(800) xor d(798) xor d(796) xor d(792) xor d(789) xor d(788) xor d(787) xor d(783) xor d(779) xor d(777) xor d(776) xor d(774) xor d(772) xor d(771) xor d(769) xor d(768) xor d(767) xor d(765) xor d(764) xor d(760) xor d(759) xor d(757) xor d(754) xor d(752) xor d(749) xor d(748) xor d(745) xor d(742) xor d(740) xor d(737) xor d(731) xor d(730) xor d(726) xor d(725) xor d(723) xor d(721) xor d(719) xor d(717) xor d(715) xor d(712) xor d(709) xor d(708) xor d(705) xor d(704) xor d(703) xor d(702) xor d(700) xor d(697) xor d(696) xor d(693) xor d(692) xor d(691) xor d(689) xor d(687) xor d(686) xor d(685) xor d(684) xor d(682) xor d(679) xor d(678) xor d(677) xor d(674) xor d(671) xor d(669) xor d(666) xor d(664) xor d(663) xor d(660) xor d(659) xor d(658) xor d(653) xor d(648) xor d(646) xor d(643) xor d(640) xor d(634) xor d(631) xor d(630) xor d(628) xor d(624) xor d(619) xor d(618) xor d(610) xor d(609) xor d(608) xor d(607) xor d(606) xor d(600) xor d(598) xor d(597) xor d(596) xor d(593) xor d(592) xor d(591) xor d(589) xor d(588) xor d(587) xor d(584) xor d(583) xor d(580) xor d(577) xor d(576) xor d(575) xor d(574) xor d(570) xor d(569) xor d(567) xor d(566) xor d(565) xor d(564) xor d(563) xor d(562) xor d(558) xor d(557) xor d(556) xor d(555) xor d(554) xor d(552) xor d(549) xor d(548) xor d(546) xor d(544) xor d(542) xor d(541) xor d(540) xor d(537) xor d(536) xor d(526) xor d(524) xor d(522) xor d(518) xor d(517) xor d(515) xor d(514) xor d(512) xor d(511) xor d(508) xor d(507) xor d(506) xor d(499) xor d(498) xor d(496) xor d(495) xor d(494) xor d(491) xor d(490) xor d(488) xor d(486) xor d(479) xor d(478) xor d(475) xor d(474) xor d(470) xor d(469) xor d(467) xor d(463) xor d(460) xor d(459) xor d(458) xor d(457) xor d(453) xor d(450) xor d(448) xor d(446) xor d(445) xor d(443) xor d(439) xor d(436) xor d(434) xor d(430) xor d(429) xor d(427) xor d(424) xor d(423) xor d(418) xor d(414) xor d(411) xor d(407) xor d(406) xor d(405) xor d(404) xor d(402) xor d(401) xor d(400) xor d(398) xor d(396) xor d(395) xor d(392) xor d(391) xor d(386) xor d(385) xor d(384) xor d(382) xor d(381) xor d(380) xor d(378) xor d(374) xor d(373) xor d(370) xor d(368) xor d(367) xor d(366) xor d(359) xor d(357) xor d(354) xor d(353) xor d(351) xor d(348) xor d(347) xor d(345) xor d(344) xor d(343) xor d(342) xor d(341) xor d(339) xor d(338) xor d(331) xor d(330) xor d(326) xor d(325) xor d(323) xor d(320) xor d(319) xor d(316) xor d(314) xor d(312) xor d(311) xor d(307) xor d(306) xor d(305) xor d(304) xor d(301) xor d(300) xor d(297) xor d(294) xor d(293) xor d(291) xor d(289) xor d(288) xor d(281) xor d(280) xor d(279) xor d(276) xor d(275) xor d(274) xor d(272) xor d(269) xor d(268) xor d(266) xor d(265) xor d(264) xor d(263) xor d(261) xor d(252) xor d(250) xor d(248) xor d(247) xor d(245) xor d(244) xor d(243) xor d(242) xor d(241) xor d(240) xor d(231) xor d(230) xor d(229) xor d(228) xor d(227) xor d(226) xor d(225) xor d(222) xor d(221) xor d(219) xor d(218) xor d(216) xor d(215) xor d(212) xor d(211) xor d(209) xor d(208) xor d(207) xor d(205) xor d(203) xor d(202) xor d(200) xor d(197) xor d(193) xor d(188) xor d(187) xor d(186) xor d(185) xor d(183) xor d(178) xor d(176) xor d(175) xor d(174) xor d(169) xor d(168) xor d(167) xor d(165) xor d(163) xor d(162) xor d(160) xor d(158) xor d(157) xor d(154) xor d(152) xor d(151) xor d(147) xor d(146) xor d(144) xor d(143) xor d(141) xor d(140) xor d(139) xor d(137) xor d(136) xor d(135) xor d(133) xor d(132) xor d(131) xor d(130) xor d(128) xor d(127) xor d(126) xor d(124) xor d(123) xor d(122) xor d(121) xor d(117) xor d(116) xor d(113) xor d(112) xor d(108) xor d(107) xor d(104) xor d(100) xor d(98) xor d(95) xor d(93) xor d(92) xor d(84) xor d(83) xor d(82) xor d(81) xor d(80) xor d(79) xor d(76) xor d(75) xor d(74) xor d(73) xor d(72) xor d(71) xor d(70) xor d(68) xor d(66) xor d(65) xor d(64) xor d(62) xor d(60) xor d(56) xor d(55) xor d(54) xor d(52) xor d(51) xor d(50) xor d(47) xor d(45) xor d(43) xor d(42) xor d(41) xor d(40) xor d(38) xor d(30) xor d(29) xor d(25) xor d(22) xor d(21) xor d(20) xor d(14) xor d(11) xor d(8) xor d(7) xor d(6) xor d(5) xor d(4) xor d(2) xor d(1) xor c(0) xor c(1) xor c(4) xor c(6) xor c(9) xor c(10) xor c(12) xor c(13) xor c(14) xor c(17) xor c(18) xor c(19) xor c(20) xor c(22) xor c(24) xor c(29) xor c(30) xor c(31);
    newcrc(7) := d(1023) xor d(1022) xor d(1021) xor d(1019) xor d(1018) xor d(1017) xor d(1016) xor d(1013) xor d(1010) xor d(1009) xor d(1008) xor d(1007) xor d(1004) xor d(1003) xor d(1002) xor d(1000) xor d(998) xor d(997) xor d(996) xor d(993) xor d(992) xor d(989) xor d(987) xor d(986) xor d(983) xor d(982) xor d(981) xor d(980) xor d(979) xor d(978) xor d(975) xor d(974) xor d(972) xor d(971) xor d(970) xor d(969) xor d(965) xor d(962) xor d(960) xor d(959) xor d(958) xor d(957) xor d(956) xor d(953) xor d(952) xor d(950) xor d(949) xor d(946) xor d(941) xor d(939) xor d(937) xor d(936) xor d(931) xor d(927) xor d(926) xor d(923) xor d(922) xor d(919) xor d(917) xor d(916) xor d(914) xor d(913) xor d(912) xor d(909) xor d(907) xor d(905) xor d(902) xor d(897) xor d(896) xor d(895) xor d(894) xor d(893) xor d(891) xor d(890) xor d(888) xor d(885) xor d(883) xor d(880) xor d(879) xor d(878) xor d(876) xor d(874) xor d(871) xor d(870) xor d(869) xor d(868) xor d(867) xor d(865) xor d(864) xor d(862) xor d(861) xor d(856) xor d(853) xor d(852) xor d(849) xor d(848) xor d(846) xor d(845) xor d(844) xor d(842) xor d(841) xor d(836) xor d(834) xor d(833) xor d(832) xor d(830) xor d(828) xor d(827) xor d(825) xor d(824) xor d(822) xor d(821) xor d(819) xor d(817) xor d(812) xor d(811) xor d(810) xor d(804) xor d(803) xor d(801) xor d(800) xor d(799) xor d(798) xor d(797) xor d(791) xor d(790) xor d(789) xor d(786) xor d(785) xor d(782) xor d(778) xor d(777) xor d(776) xor d(775) xor d(774) xor d(773) xor d(772) xor d(770) xor d(768) xor d(767) xor d(766) xor d(763) xor d(762) xor d(761) xor d(760) xor d(756) xor d(749) xor d(748) xor d(747) xor d(746) xor d(744) xor d(743) xor d(742) xor d(740) xor d(738) xor d(736) xor d(729) xor d(726) xor d(725) xor d(723) xor d(721) xor d(719) xor d(718) xor d(716) xor d(715) xor d(713) xor d(709) xor d(708) xor d(707) xor d(706) xor d(705) xor d(703) xor d(702) xor d(700) xor d(697) xor d(695) xor d(692) xor d(691) xor d(690) xor d(689) xor d(688) xor d(685) xor d(683) xor d(679) xor d(678) xor d(674) xor d(673) xor d(669) xor d(668) xor d(666) xor d(664) xor d(661) xor d(660) xor d(659) xor d(658) xor d(656) xor d(655) xor d(654) xor d(653) xor d(652) xor d(648) xor d(647) xor d(646) xor d(642) xor d(641) xor d(640) xor d(636) xor d(635) xor d(631) xor d(630) xor d(626) xor d(625) xor d(624) xor d(623) xor d(617) xor d(615) xor d(613) xor d(612) xor d(608) xor d(606) xor d(604) xor d(603) xor d(602) xor d(601) xor d(600) xor d(598) xor d(597) xor d(596) xor d(595) xor d(594) xor d(591) xor d(590) xor d(589) xor d(588) xor d(587) xor d(586) xor d(584) xor d(583) xor d(581) xor d(580) xor d(577) xor d(576) xor d(574) xor d(573) xor d(570) xor d(568) xor d(566) xor d(564) xor d(561) xor d(560) xor d(559) xor d(554) xor d(553) xor d(551) xor d(550) xor d(547) xor d(543) xor d(541) xor d(540) xor d(539) xor d(538) xor d(537) xor d(535) xor d(534) xor d(532) xor d(531) xor d(530) xor d(529) xor d(528) xor d(527) xor d(526) xor d(523) xor d(522) xor d(521) xor d(515) xor d(514) xor d(513) xor d(511) xor d(510) xor d(509) xor d(506) xor d(502) xor d(501) xor d(499) xor d(497) xor d(496) xor d(494) xor d(493) xor d(490) xor d(488) xor d(487) xor d(486) xor d(483) xor d(482) xor d(481) xor d(477) xor d(475) xor d(472) xor d(471) xor d(465) xor d(462) xor d(460) xor d(459) xor d(454) xor d(452) xor d(451) xor d(450) xor d(448) xor d(447) xor d(446) xor d(440) xor d(436) xor d(435) xor d(434) xor d(433) xor d(431) xor d(430) xor d(428) xor d(425) xor d(422) xor d(418) xor d(416) xor d(415) xor d(414) xor d(409) xor d(406) xor d(404) xor d(403) xor d(402) xor d(401) xor d(400) xor d(398) xor d(397) xor d(391) xor d(390) xor d(388) xor d(385) xor d(383) xor d(382) xor d(379) xor d(378) xor d(376) xor d(375) xor d(372) xor d(371) xor d(367) xor d(366) xor d(363) xor d(362) xor d(360) xor d(359) xor d(357) xor d(355) xor d(354) xor d(353) xor d(352) xor d(347) xor d(346) xor d(343) xor d(341) xor d(340) xor d(338) xor d(337) xor d(335) xor d(334) xor d(333) xor d(332) xor d(331) xor d(328) xor d(326) xor d(324) xor d(322) xor d(319) xor d(318) xor d(313) xor d(310) xor d(309) xor d(308) xor d(307) xor d(306) xor d(303) xor d(301) xor d(300) xor d(299) xor d(297) xor d(296) xor d(289) xor d(288) xor d(287) xor d(286) xor d(283) xor d(282) xor d(281) xor d(280) xor d(279) xor d(275) xor d(274) xor d(270) xor d(268) xor d(267) xor d(266) xor d(262) xor d(261) xor d(259) xor d(257) xor d(255) xor d(253) xor d(252) xor d(251) xor d(249) xor d(246) xor d(245) xor d(244) xor d(242) xor d(241) xor d(237) xor d(234) xor d(232) xor d(231) xor d(229) xor d(224) xor d(223) xor d(222) xor d(220) xor d(219) xor d(217) xor d(214) xor d(213) xor d(207) xor d(206) xor d(204) xor d(202) xor d(199) xor d(197) xor d(193) xor d(192) xor d(191) xor d(190) xor d(189) xor d(187) xor d(184) xor d(183) xor d(182) xor d(179) xor d(177) xor d(176) xor d(175) xor d(172) xor d(171) xor d(168) xor d(167) xor d(164) xor d(163) xor d(162) xor d(159) xor d(156) xor d(153) xor d(152) xor d(151) xor d(149) xor d(148) xor d(147) xor d(145) xor d(143) xor d(142) xor d(141) xor d(140) xor d(138) xor d(135) xor d(133) xor d(131) xor d(129) xor d(126) xor d(124) xor d(122) xor d(119) xor d(116) xor d(111) xor d(110) xor d(109) xor d(108) xor d(106) xor d(105) xor d(104) xor d(103) xor d(98) xor d(97) xor d(95) xor d(93) xor d(87) xor d(80) xor d(79) xor d(77) xor d(76) xor d(75) xor d(74) xor d(71) xor d(69) xor d(68) xor d(60) xor d(58) xor d(57) xor d(56) xor d(54) xor d(52) xor d(51) xor d(50) xor d(47) xor d(46) xor d(45) xor d(43) xor d(42) xor d(41) xor d(39) xor d(37) xor d(34) xor d(32) xor d(29) xor d(28) xor d(25) xor d(24) xor d(23) xor d(22) xor d(21) xor d(16) xor d(15) xor d(10) xor d(8) xor d(7) xor d(5) xor d(3) xor d(2) xor d(0) xor c(0) xor c(1) xor c(4) xor c(5) xor c(6) xor c(8) xor c(10) xor c(11) xor c(12) xor c(15) xor c(16) xor c(17) xor c(18) xor c(21) xor c(24) xor c(25) xor c(26) xor c(27) xor c(29) xor c(30) xor c(31);
    newcrc(8) := d(1023) xor d(1022) xor d(1021) xor d(1020) xor d(1017) xor d(1016) xor d(1015) xor d(1014) xor d(1012) xor d(1010) xor d(1006) xor d(1003) xor d(1001) xor d(1000) xor d(997) xor d(996) xor d(993) xor d(992) xor d(988) xor d(987) xor d(985) xor d(978) xor d(977) xor d(976) xor d(974) xor d(973) xor d(972) xor d(970) xor d(967) xor d(966) xor d(963) xor d(961) xor d(957) xor d(955) xor d(951) xor d(948) xor d(947) xor d(944) xor d(942) xor d(941) xor d(940) xor d(939) xor d(937) xor d(935) xor d(934) xor d(933) xor d(932) xor d(931) xor d(928) xor d(927) xor d(924) xor d(923) xor d(914) xor d(913) xor d(908) xor d(907) xor d(904) xor d(902) xor d(901) xor d(900) xor d(899) xor d(895) xor d(894) xor d(893) xor d(892) xor d(890) xor d(887) xor d(884) xor d(883) xor d(880) xor d(878) xor d(876) xor d(874) xor d(873) xor d(872) xor d(870) xor d(867) xor d(866) xor d(865) xor d(862) xor d(861) xor d(860) xor d(859) xor d(851) xor d(848) xor d(847) xor d(845) xor d(843) xor d(840) xor d(839) xor d(833) xor d(832) xor d(831) xor d(829) xor d(828) xor d(827) xor d(826) xor d(824) xor d(823) xor d(822) xor d(820) xor d(819) xor d(816) xor d(815) xor d(814) xor d(810) xor d(809) xor d(808) xor d(807) xor d(806) xor d(805) xor d(803) xor d(801) xor d(799) xor d(793) xor d(792) xor d(790) xor d(788) xor d(787) xor d(785) xor d(784) xor d(783) xor d(782) xor d(780) xor d(779) xor d(778) xor d(777) xor d(775) xor d(773) xor d(771) xor d(768) xor d(765) xor d(764) xor d(761) xor d(758) xor d(757) xor d(756) xor d(755) xor d(753) xor d(749) xor d(745) xor d(743) xor d(742) xor d(740) xor d(739) xor d(737) xor d(736) xor d(732) xor d(731) xor d(730) xor d(729) xor d(726) xor d(725) xor d(723) xor d(721) xor d(717) xor d(716) xor d(715) xor d(714) xor d(709) xor d(706) xor d(703) xor d(702) xor d(700) xor d(696) xor d(695) xor d(694) xor d(692) xor d(690) xor d(687) xor d(684) xor d(679) xor d(673) xor d(672) xor d(668) xor d(666) xor d(662) xor d(661) xor d(660) xor d(659) xor d(658) xor d(657) xor d(654) xor d(652) xor d(647) xor d(646) xor d(644) xor d(643) xor d(641) xor d(640) xor d(637) xor d(631) xor d(630) xor d(629) xor d(627) xor d(625) xor d(623) xor d(620) xor d(619) xor d(618) xor d(617) xor d(616) xor d(615) xor d(614) xor d(612) xor d(611) xor d(610) xor d(606) xor d(605) xor d(601) xor d(600) xor d(598) xor d(597) xor d(593) xor d(590) xor d(589) xor d(588) xor d(586) xor d(584) xor d(583) xor d(582) xor d(581) xor d(580) xor d(577) xor d(573) xor d(569) xor d(563) xor d(562) xor d(558) xor d(557) xor d(556) xor d(552) xor d(549) xor d(548) xor d(545) xor d(544) xor d(541) xor d(538) xor d(536) xor d(534) xor d(533) xor d(527) xor d(526) xor d(525) xor d(524) xor d(523) xor d(521) xor d(519) xor d(518) xor d(515) xor d(508) xor d(506) xor d(503) xor d(501) xor d(498) xor d(497) xor d(493) xor d(492) xor d(490) xor d(487) xor d(486) xor d(484) xor d(481) xor d(480) xor d(479) xor d(478) xor d(477) xor d(473) xor d(470) xor d(468) xor d(466) xor d(465) xor d(464) xor d(463) xor d(462) xor d(460) xor d(458) xor d(455) xor d(453) xor d(451) xor d(450) xor d(447) xor d(444) xor d(441) xor d(435) xor d(433) xor d(432) xor d(431) xor d(429) xor d(426) xor d(424) xor d(423) xor d(422) xor d(418) xor d(417) xor d(415) xor d(414) xor d(412) xor d(410) xor d(409) xor d(408) xor d(403) xor d(402) xor d(401) xor d(400) xor d(396) xor d(393) xor d(390) xor d(389) xor d(388) xor d(387) xor d(384) xor d(383) xor d(381) xor d(380) xor d(379) xor d(378) xor d(377) xor d(374) xor d(373) xor d(369) xor d(367) xor d(366) xor d(364) xor d(362) xor d(361) xor d(360) xor d(359) xor d(357) xor d(356) xor d(355) xor d(354) xor d(349) xor d(345) xor d(337) xor d(336) xor d(332) xor d(329) xor d(328) xor d(325) xor d(323) xor d(322) xor d(321) xor d(318) xor d(317) xor d(315) xor d(314) xor d(312) xor d(311) xor d(308) xor d(307) xor d(305) xor d(304) xor d(303) xor d(301) xor d(299) xor d(296) xor d(295) xor d(294) xor d(292) xor d(289) xor d(286) xor d(284) xor d(282) xor d(281) xor d(280) xor d(279) xor d(277) xor d(275) xor d(274) xor d(273) xor d(271) xor d(267) xor d(265) xor d(264) xor d(263) xor d(262) xor d(261) xor d(260) xor d(259) xor d(258) xor d(257) xor d(256) xor d(255) xor d(254) xor d(253) xor d(250) xor d(248) xor d(247) xor d(246) xor d(245) xor d(242) xor d(238) xor d(237) xor d(235) xor d(234) xor d(233) xor d(232) xor d(228) xor d(227) xor d(226) xor d(225) xor d(223) xor d(221) xor d(220) xor d(218) xor d(216) xor d(215) xor d(212) xor d(210) xor d(209) xor d(205) xor d(202) xor d(201) xor d(200) xor d(199) xor d(197) xor d(186) xor d(185) xor d(184) xor d(182) xor d(180) xor d(178) xor d(177) xor d(176) xor d(173) xor d(171) xor d(170) xor d(168) xor d(167) xor d(166) xor d(165) xor d(164) xor d(163) xor d(162) xor d(161) xor d(160) xor d(158) xor d(157) xor d(156) xor d(155) xor d(154) xor d(153) xor d(152) xor d(151) xor d(150) xor d(148) xor d(146) xor d(142) xor d(141) xor d(139) xor d(137) xor d(135) xor d(130) xor d(128) xor d(126) xor d(120) xor d(119) xor d(118) xor d(116) xor d(114) xor d(113) xor d(112) xor d(109) xor d(107) xor d(105) xor d(103) xor d(101) xor d(97) xor d(95) xor d(88) xor d(87) xor d(85) xor d(84) xor d(83) xor d(82) xor d(80) xor d(79) xor d(78) xor d(77) xor d(76) xor d(75) xor d(73) xor d(70) xor d(69) xor d(68) xor d(67) xor d(66) xor d(65) xor d(63) xor d(60) xor d(59) xor d(57) xor d(54) xor d(52) xor d(51) xor d(50) xor d(46) xor d(45) xor d(43) xor d(42) xor d(40) xor d(38) xor d(37) xor d(35) xor d(34) xor d(33) xor d(32) xor d(31) xor d(28) xor d(23) xor d(22) xor d(17) xor d(12) xor d(11) xor d(10) xor d(8) xor d(4) xor d(3) xor d(1) xor d(0) xor c(0) xor c(1) xor c(4) xor c(5) xor c(8) xor c(9) xor c(11) xor c(14) xor c(18) xor c(20) xor c(22) xor c(23) xor c(24) xor c(25) xor c(28) xor c(29) xor c(30) xor c(31);
    newcrc(9) := d(1023) xor d(1022) xor d(1021) xor d(1018) xor d(1017) xor d(1016) xor d(1015) xor d(1013) xor d(1011) xor d(1007) xor d(1004) xor d(1002) xor d(1001) xor d(998) xor d(997) xor d(994) xor d(993) xor d(989) xor d(988) xor d(986) xor d(979) xor d(978) xor d(977) xor d(975) xor d(974) xor d(973) xor d(971) xor d(968) xor d(967) xor d(964) xor d(962) xor d(958) xor d(956) xor d(952) xor d(949) xor d(948) xor d(945) xor d(943) xor d(942) xor d(941) xor d(940) xor d(938) xor d(936) xor d(935) xor d(934) xor d(933) xor d(932) xor d(929) xor d(928) xor d(925) xor d(924) xor d(915) xor d(914) xor d(909) xor d(908) xor d(905) xor d(903) xor d(902) xor d(901) xor d(900) xor d(896) xor d(895) xor d(894) xor d(893) xor d(891) xor d(888) xor d(885) xor d(884) xor d(881) xor d(879) xor d(877) xor d(875) xor d(874) xor d(873) xor d(871) xor d(868) xor d(867) xor d(866) xor d(863) xor d(862) xor d(861) xor d(860) xor d(852) xor d(849) xor d(848) xor d(846) xor d(844) xor d(841) xor d(840) xor d(834) xor d(833) xor d(832) xor d(830) xor d(829) xor d(828) xor d(827) xor d(825) xor d(824) xor d(823) xor d(821) xor d(820) xor d(817) xor d(816) xor d(815) xor d(811) xor d(810) xor d(809) xor d(808) xor d(807) xor d(806) xor d(804) xor d(802) xor d(800) xor d(794) xor d(793) xor d(791) xor d(789) xor d(788) xor d(786) xor d(785) xor d(784) xor d(783) xor d(781) xor d(780) xor d(779) xor d(778) xor d(776) xor d(774) xor d(772) xor d(769) xor d(766) xor d(765) xor d(762) xor d(759) xor d(758) xor d(757) xor d(756) xor d(754) xor d(750) xor d(746) xor d(744) xor d(743) xor d(741) xor d(740) xor d(738) xor d(737) xor d(733) xor d(732) xor d(731) xor d(730) xor d(727) xor d(726) xor d(724) xor d(722) xor d(718) xor d(717) xor d(716) xor d(715) xor d(710) xor d(707) xor d(704) xor d(703) xor d(701) xor d(697) xor d(696) xor d(695) xor d(693) xor d(691) xor d(688) xor d(685) xor d(680) xor d(674) xor d(673) xor d(669) xor d(667) xor d(663) xor d(662) xor d(661) xor d(660) xor d(659) xor d(658) xor d(655) xor d(653) xor d(648) xor d(647) xor d(645) xor d(644) xor d(642) xor d(641) xor d(638) xor d(632) xor d(631) xor d(630) xor d(628) xor d(626) xor d(624) xor d(621) xor d(620) xor d(619) xor d(618) xor d(617) xor d(616) xor d(615) xor d(613) xor d(612) xor d(611) xor d(607) xor d(606) xor d(602) xor d(601) xor d(599) xor d(598) xor d(594) xor d(591) xor d(590) xor d(589) xor d(587) xor d(585) xor d(584) xor d(583) xor d(582) xor d(581) xor d(578) xor d(574) xor d(570) xor d(564) xor d(563) xor d(559) xor d(558) xor d(557) xor d(553) xor d(550) xor d(549) xor d(546) xor d(545) xor d(542) xor d(539) xor d(537) xor d(535) xor d(534) xor d(528) xor d(527) xor d(526) xor d(525) xor d(524) xor d(522) xor d(520) xor d(519) xor d(516) xor d(509) xor d(507) xor d(504) xor d(502) xor d(499) xor d(498) xor d(494) xor d(493) xor d(491) xor d(488) xor d(487) xor d(485) xor d(482) xor d(481) xor d(480) xor d(479) xor d(478) xor d(474) xor d(471) xor d(469) xor d(467) xor d(466) xor d(465) xor d(464) xor d(463) xor d(461) xor d(459) xor d(456) xor d(454) xor d(452) xor d(451) xor d(448) xor d(445) xor d(442) xor d(436) xor d(434) xor d(433) xor d(432) xor d(430) xor d(427) xor d(425) xor d(424) xor d(423) xor d(419) xor d(418) xor d(416) xor d(415) xor d(413) xor d(411) xor d(410) xor d(409) xor d(404) xor d(403) xor d(402) xor d(401) xor d(397) xor d(394) xor d(391) xor d(390) xor d(389) xor d(388) xor d(385) xor d(384) xor d(382) xor d(381) xor d(380) xor d(379) xor d(378) xor d(375) xor d(374) xor d(370) xor d(368) xor d(367) xor d(365) xor d(363) xor d(362) xor d(361) xor d(360) xor d(358) xor d(357) xor d(356) xor d(355) xor d(350) xor d(346) xor d(338) xor d(337) xor d(333) xor d(330) xor d(329) xor d(326) xor d(324) xor d(323) xor d(322) xor d(319) xor d(318) xor d(316) xor d(315) xor d(313) xor d(312) xor d(309) xor d(308) xor d(306) xor d(305) xor d(304) xor d(302) xor d(300) xor d(297) xor d(296) xor d(295) xor d(293) xor d(290) xor d(287) xor d(285) xor d(283) xor d(282) xor d(281) xor d(280) xor d(278) xor d(276) xor d(275) xor d(274) xor d(272) xor d(268) xor d(266) xor d(265) xor d(264) xor d(263) xor d(262) xor d(261) xor d(260) xor d(259) xor d(258) xor d(257) xor d(256) xor d(255) xor d(254) xor d(251) xor d(249) xor d(248) xor d(247) xor d(246) xor d(243) xor d(239) xor d(238) xor d(236) xor d(235) xor d(234) xor d(233) xor d(229) xor d(228) xor d(227) xor d(226) xor d(224) xor d(222) xor d(221) xor d(219) xor d(217) xor d(216) xor d(213) xor d(211) xor d(210) xor d(206) xor d(203) xor d(202) xor d(201) xor d(200) xor d(198) xor d(187) xor d(186) xor d(185) xor d(183) xor d(181) xor d(179) xor d(178) xor d(177) xor d(174) xor d(172) xor d(171) xor d(169) xor d(168) xor d(167) xor d(166) xor d(165) xor d(164) xor d(163) xor d(162) xor d(161) xor d(159) xor d(158) xor d(157) xor d(156) xor d(155) xor d(154) xor d(153) xor d(152) xor d(151) xor d(149) xor d(147) xor d(143) xor d(142) xor d(140) xor d(138) xor d(136) xor d(131) xor d(129) xor d(127) xor d(121) xor d(120) xor d(119) xor d(117) xor d(115) xor d(114) xor d(113) xor d(110) xor d(108) xor d(106) xor d(104) xor d(102) xor d(98) xor d(96) xor d(89) xor d(88) xor d(86) xor d(85) xor d(84) xor d(83) xor d(81) xor d(80) xor d(79) xor d(78) xor d(77) xor d(76) xor d(74) xor d(71) xor d(70) xor d(69) xor d(68) xor d(67) xor d(66) xor d(64) xor d(61) xor d(60) xor d(58) xor d(55) xor d(53) xor d(52) xor d(51) xor d(47) xor d(46) xor d(44) xor d(43) xor d(41) xor d(39) xor d(38) xor d(36) xor d(35) xor d(34) xor d(33) xor d(32) xor d(29) xor d(24) xor d(23) xor d(18) xor d(13) xor d(12) xor d(11) xor d(9) xor d(5) xor d(4) xor d(2) xor d(1) xor c(1) xor c(2) xor c(5) xor c(6) xor c(9) xor c(10) xor c(12) xor c(15) xor c(19) xor c(21) xor c(23) xor c(24) xor c(25) xor c(26) xor c(29) xor c(30) xor c(31);
    newcrc(10) := d(1023) xor d(1022) xor d(1021) xor d(1017) xor d(1015) xor d(1014) xor d(1011) xor d(1009) xor d(1006) xor d(1004) xor d(1003) xor d(1002) xor d(1000) xor d(996) xor d(995) xor d(992) xor d(989) xor d(987) xor d(985) xor d(984) xor d(983) xor d(982) xor d(981) xor d(977) xor d(976) xor d(972) xor d(971) xor d(969) xor d(968) xor d(967) xor d(965) xor d(963) xor d(960) xor d(958) xor d(957) xor d(955) xor d(954) xor d(949) xor d(948) xor d(946) xor d(943) xor d(942) xor d(938) xor d(937) xor d(936) xor d(931) xor d(930) xor d(929) xor d(926) xor d(925) xor d(920) xor d(918) xor d(917) xor d(916) xor d(909) xor d(907) xor d(900) xor d(899) xor d(898) xor d(895) xor d(894) xor d(893) xor d(892) xor d(891) xor d(890) xor d(887) xor d(885) xor d(883) xor d(882) xor d(881) xor d(880) xor d(879) xor d(877) xor d(873) xor d(872) xor d(871) xor d(864) xor d(862) xor d(860) xor d(859) xor d(857) xor d(854) xor d(851) xor d(848) xor d(847) xor d(846) xor d(845) xor d(841) xor d(840) xor d(839) xor d(837) xor d(833) xor d(832) xor d(831) xor d(830) xor d(829) xor d(828) xor d(827) xor d(826) xor d(822) xor d(821) xor d(819) xor d(817) xor d(815) xor d(814) xor d(813) xor d(806) xor d(805) xor d(804) xor d(802) xor d(801) xor d(800) xor d(798) xor d(795) xor d(794) xor d(793) xor d(792) xor d(791) xor d(790) xor d(789) xor d(788) xor d(787) xor d(781) xor d(779) xor d(777) xor d(776) xor d(775) xor d(774) xor d(773) xor d(770) xor d(769) xor d(766) xor d(765) xor d(762) xor d(760) xor d(759) xor d(757) xor d(756) xor d(753) xor d(751) xor d(750) xor d(748) xor d(745) xor d(740) xor d(739) xor d(738) xor d(736) xor d(734) xor d(733) xor d(729) xor d(728) xor d(724) xor d(722) xor d(721) xor d(720) xor d(718) xor d(717) xor d(716) xor d(715) xor d(711) xor d(710) xor d(707) xor d(705) xor d(701) xor d(700) xor d(697) xor d(696) xor d(695) xor d(693) xor d(692) xor d(691) xor d(687) xor d(681) xor d(680) xor d(673) xor d(672) xor d(669) xor d(667) xor d(666) xor d(665) xor d(664) xor d(663) xor d(662) xor d(661) xor d(660) xor d(659) xor d(658) xor d(655) xor d(654) xor d(653) xor d(652) xor d(645) xor d(644) xor d(643) xor d(640) xor d(639) xor d(636) xor d(633) xor d(631) xor d(630) xor d(627) xor d(626) xor d(625) xor d(624) xor d(623) xor d(622) xor d(621) xor d(618) xor d(616) xor d(615) xor d(614) xor d(611) xor d(610) xor d(609) xor d(608) xor d(606) xor d(604) xor d(596) xor d(593) xor d(590) xor d(588) xor d(587) xor d(584) xor d(582) xor d(580) xor d(579) xor d(578) xor d(574) xor d(573) xor d(567) xor d(564) xor d(563) xor d(561) xor d(559) xor d(557) xor d(556) xor d(555) xor d(550) xor d(549) xor d(547) xor d(546) xor d(545) xor d(543) xor d(542) xor d(539) xor d(538) xor d(536) xor d(534) xor d(532) xor d(531) xor d(530) xor d(527) xor d(523) xor d(522) xor d(520) xor d(519) xor d(518) xor d(517) xor d(516) xor d(514) xor d(512) xor d(511) xor d(507) xor d(506) xor d(505) xor d(503) xor d(502) xor d(501) xor d(499) xor d(493) xor d(491) xor d(490) xor d(477) xor d(476) xor d(475) xor d(467) xor d(466) xor d(461) xor d(460) xor d(458) xor d(457) xor d(455) xor d(453) xor d(450) xor d(448) xor d(446) xor d(444) xor d(443) xor d(436) xor d(435) xor d(431) xor d(428) xor d(426) xor d(425) xor d(422) xor d(420) xor d(418) xor d(417) xor d(411) xor d(410) xor d(409) xor d(408) xor d(407) xor d(403) xor d(402) xor d(400) xor d(399) xor d(396) xor d(395) xor d(393) xor d(389) xor d(388) xor d(387) xor d(385) xor d(383) xor d(382) xor d(380) xor d(379) xor d(378) xor d(375) xor d(374) xor d(372) xor d(371) xor d(364) xor d(361) xor d(356) xor d(353) xor d(351) xor d(349) xor d(348) xor d(345) xor d(344) xor d(342) xor d(341) xor d(337) xor d(335) xor d(333) xor d(331) xor d(330) xor d(328) xor d(325) xor d(324) xor d(323) xor d(322) xor d(321) xor d(318) xor d(316) xor d(315) xor d(314) xor d(313) xor d(312) xor d(307) xor d(306) xor d(302) xor d(301) xor d(300) xor d(299) xor d(295) xor d(292) xor d(291) xor d(290) xor d(287) xor d(284) xor d(282) xor d(281) xor d(275) xor d(274) xor d(268) xor d(267) xor d(266) xor d(263) xor d(262) xor d(260) xor d(258) xor d(256) xor d(250) xor d(249) xor d(247) xor d(244) xor d(243) xor d(240) xor d(239) xor d(236) xor d(235) xor d(229) xor d(226) xor d(225) xor d(224) xor d(223) xor d(222) xor d(220) xor d(218) xor d(217) xor d(216) xor d(211) xor d(210) xor d(209) xor d(208) xor d(204) xor d(198) xor d(197) xor d(194) xor d(193) xor d(192) xor d(191) xor d(190) xor d(187) xor d(184) xor d(183) xor d(180) xor d(179) xor d(178) xor d(175) xor d(173) xor d(171) xor d(168) xor d(165) xor d(164) xor d(163) xor d(161) xor d(160) xor d(159) xor d(157) xor d(154) xor d(153) xor d(152) xor d(151) xor d(150) xor d(149) xor d(148) xor d(141) xor d(139) xor d(136) xor d(135) xor d(134) xor d(130) xor d(127) xor d(126) xor d(125) xor d(123) xor d(122) xor d(121) xor d(120) xor d(119) xor d(117) xor d(115) xor d(113) xor d(110) xor d(109) xor d(107) xor d(106) xor d(105) xor d(104) xor d(101) xor d(98) xor d(96) xor d(95) xor d(94) xor d(90) xor d(89) xor d(86) xor d(83) xor d(80) xor d(78) xor d(77) xor d(75) xor d(73) xor d(71) xor d(70) xor d(69) xor d(66) xor d(63) xor d(62) xor d(60) xor d(59) xor d(58) xor d(56) xor d(55) xor d(52) xor d(50) xor d(42) xor d(40) xor d(39) xor d(36) xor d(35) xor d(33) xor d(32) xor d(31) xor d(29) xor d(28) xor d(26) xor d(19) xor d(16) xor d(14) xor d(13) xor d(9) xor d(5) xor d(3) xor d(2) xor d(0) xor c(0) xor c(3) xor c(4) xor c(8) xor c(10) xor c(11) xor c(12) xor c(14) xor c(17) xor c(19) xor c(22) xor c(23) xor c(25) xor c(29) xor c(30) xor c(31);
    newcrc(11) := d(1023) xor d(1022) xor d(1021) xor d(1019) xor d(1011) xor d(1010) xor d(1009) xor d(1008) xor d(1007) xor d(1006) xor d(1003) xor d(1001) xor d(1000) xor d(999) xor d(998) xor d(997) xor d(994) xor d(993) xor d(992) xor d(988) xor d(986) xor d(981) xor d(980) xor d(979) xor d(975) xor d(974) xor d(973) xor d(972) xor d(971) xor d(970) xor d(969) xor d(968) xor d(967) xor d(966) xor d(964) xor d(961) xor d(960) xor d(956) xor d(954) xor d(953) xor d(949) xor d(948) xor d(947) xor d(943) xor d(941) xor d(937) xor d(935) xor d(934) xor d(933) xor d(932) xor d(930) xor d(927) xor d(926) xor d(921) xor d(920) xor d(919) xor d(915) xor d(908) xor d(907) xor d(906) xor d(904) xor d(903) xor d(902) xor d(898) xor d(897) xor d(895) xor d(894) xor d(892) xor d(890) xor d(889) xor d(888) xor d(887) xor d(884) xor d(882) xor d(880) xor d(879) xor d(877) xor d(876) xor d(875) xor d(872) xor d(871) xor d(869) xor d(868) xor d(867) xor d(865) xor d(859) xor d(858) xor d(857) xor d(855) xor d(854) xor d(853) xor d(852) xor d(851) xor d(850) xor d(847) xor d(841) xor d(839) xor d(838) xor d(837) xor d(835) xor d(833) xor d(831) xor d(830) xor d(829) xor d(828) xor d(825) xor d(824) xor d(823) xor d(822) xor d(820) xor d(819) xor d(813) xor d(812) xor d(811) xor d(810) xor d(809) xor d(808) xor d(805) xor d(804) xor d(801) xor d(800) xor d(799) xor d(798) xor d(796) xor d(795) xor d(794) xor d(792) xor d(790) xor d(789) xor d(786) xor d(785) xor d(784) xor d(778) xor d(777) xor d(775) xor d(771) xor d(770) xor d(769) xor d(766) xor d(765) xor d(762) xor d(761) xor d(760) xor d(757) xor d(756) xor d(755) xor d(754) xor d(753) xor d(752) xor d(751) xor d(750) xor d(749) xor d(748) xor d(747) xor d(746) xor d(744) xor d(742) xor d(739) xor d(737) xor d(736) xor d(735) xor d(734) xor d(732) xor d(731) xor d(730) xor d(727) xor d(724) xor d(720) xor d(718) xor d(717) xor d(716) xor d(715) xor d(712) xor d(711) xor d(710) xor d(707) xor d(706) xor d(704) xor d(700) xor d(697) xor d(696) xor d(695) xor d(692) xor d(691) xor d(689) xor d(688) xor d(687) xor d(686) xor d(682) xor d(681) xor d(680) xor d(675) xor d(672) xor d(669) xor d(664) xor d(663) xor d(662) xor d(661) xor d(660) xor d(659) xor d(658) xor d(654) xor d(652) xor d(649) xor d(648) xor d(645) xor d(642) xor d(641) xor d(637) xor d(636) xor d(634) xor d(631) xor d(630) xor d(629) xor d(628) xor d(627) xor d(625) xor d(622) xor d(620) xor d(616) xor d(613) xor d(606) xor d(605) xor d(604) xor d(603) xor d(602) xor d(600) xor d(599) xor d(597) xor d(596) xor d(595) xor d(594) xor d(593) xor d(592) xor d(589) xor d(588) xor d(587) xor d(586) xor d(581) xor d(579) xor d(578) xor d(573) xor d(571) xor d(568) xor d(567) xor d(564) xor d(563) xor d(562) xor d(561) xor d(555) xor d(554) xor d(550) xor d(549) xor d(548) xor d(547) xor d(546) xor d(545) xor d(544) xor d(543) xor d(542) xor d(537) xor d(534) xor d(533) xor d(530) xor d(529) xor d(526) xor d(525) xor d(524) xor d(523) xor d(522) xor d(520) xor d(517) xor d(516) xor d(515) xor d(514) xor d(513) xor d(511) xor d(510) xor d(504) xor d(503) xor d(501) xor d(495) xor d(493) xor d(490) xor d(489) xor d(488) xor d(486) xor d(483) xor d(482) xor d(481) xor d(480) xor d(479) xor d(478) xor d(472) xor d(470) xor d(467) xor d(465) xor d(464) xor d(459) xor d(456) xor d(454) xor d(452) xor d(451) xor d(450) xor d(448) xor d(447) xor d(445) xor d(434) xor d(433) xor d(432) xor d(429) xor d(427) xor d(426) xor d(424) xor d(423) xor d(422) xor d(421) xor d(416) xor d(414) xor d(411) xor d(410) xor d(407) xor d(405) xor d(403) xor d(401) xor d(399) xor d(398) xor d(397) xor d(394) xor d(393) xor d(392) xor d(391) xor d(389) xor d(387) xor d(384) xor d(383) xor d(380) xor d(379) xor d(378) xor d(375) xor d(374) xor d(373) xor d(369) xor d(368) xor d(366) xor d(365) xor d(363) xor d(359) xor d(358) xor d(354) xor d(353) xor d(352) xor d(350) xor d(348) xor d(347) xor d(346) xor d(344) xor d(343) xor d(341) xor d(339) xor d(337) xor d(336) xor d(335) xor d(333) xor d(332) xor d(331) xor d(329) xor d(328) xor d(327) xor d(326) xor d(325) xor d(324) xor d(323) xor d(321) xor d(320) xor d(318) xor d(316) xor d(314) xor d(313) xor d(312) xor d(310) xor d(309) xor d(308) xor d(307) xor d(305) xor d(301) xor d(299) xor d(298) xor d(297) xor d(295) xor d(294) xor d(293) xor d(291) xor d(290) xor d(287) xor d(286) xor d(285) xor d(282) xor d(279) xor d(277) xor d(275) xor d(274) xor d(273) xor d(267) xor d(265) xor d(263) xor d(255) xor d(252) xor d(251) xor d(250) xor d(245) xor d(244) xor d(243) xor d(241) xor d(240) xor d(236) xor d(234) xor d(228) xor d(225) xor d(223) xor d(221) xor d(219) xor d(218) xor d(217) xor d(216) xor d(214) xor d(211) xor d(208) xor d(207) xor d(205) xor d(203) xor d(202) xor d(201) xor d(197) xor d(195) xor d(190) xor d(186) xor d(185) xor d(184) xor d(183) xor d(182) xor d(181) xor d(180) xor d(179) xor d(176) xor d(174) xor d(171) xor d(170) xor d(167) xor d(165) xor d(164) xor d(160) xor d(156) xor d(154) xor d(153) xor d(152) xor d(150) xor d(144) xor d(143) xor d(142) xor d(140) xor d(134) xor d(132) xor d(131) xor d(125) xor d(124) xor d(122) xor d(121) xor d(120) xor d(119) xor d(117) xor d(113) xor d(108) xor d(107) xor d(105) xor d(104) xor d(103) xor d(102) xor d(101) xor d(98) xor d(94) xor d(91) xor d(90) xor d(85) xor d(83) xor d(82) xor d(78) xor d(76) xor d(74) xor d(73) xor d(71) xor d(70) xor d(68) xor d(66) xor d(65) xor d(64) xor d(59) xor d(58) xor d(57) xor d(56) xor d(55) xor d(54) xor d(51) xor d(50) xor d(48) xor d(47) xor d(45) xor d(44) xor d(43) xor d(41) xor d(40) xor d(36) xor d(33) xor d(31) xor d(28) xor d(27) xor d(26) xor d(25) xor d(24) xor d(20) xor d(17) xor d(16) xor d(15) xor d(14) xor d(12) xor d(9) xor d(4) xor d(3) xor d(1) xor d(0) xor c(0) xor c(1) xor c(2) xor c(5) xor c(6) xor c(7) xor c(8) xor c(9) xor c(11) xor c(14) xor c(15) xor c(16) xor c(17) xor c(18) xor c(19) xor c(27) xor c(29) xor c(30) xor c(31);
    newcrc(12) := d(1023) xor d(1022) xor d(1021) xor d(1020) xor d(1019) xor d(1018) xor d(1016) xor d(1015) xor d(1010) xor d(1007) xor d(1006) xor d(1005) xor d(1002) xor d(1001) xor d(996) xor d(995) xor d(993) xor d(992) xor d(990) xor d(989) xor d(987) xor d(985) xor d(984) xor d(983) xor d(979) xor d(978) xor d(977) xor d(976) xor d(973) xor d(972) xor d(970) xor d(969) xor d(968) xor d(965) xor d(962) xor d(961) xor d(960) xor d(959) xor d(958) xor d(957) xor d(953) xor d(949) xor d(942) xor d(941) xor d(939) xor d(936) xor d(928) xor d(927) xor d(922) xor d(921) xor d(918) xor d(917) xor d(916) xor d(915) xor d(910) xor d(909) xor d(908) xor d(906) xor d(905) xor d(902) xor d(901) xor d(900) xor d(897) xor d(895) xor d(888) xor d(887) xor d(886) xor d(885) xor d(880) xor d(879) xor d(875) xor d(874) xor d(872) xor d(871) xor d(870) xor d(867) xor d(866) xor d(863) xor d(861) xor d(858) xor d(857) xor d(856) xor d(855) xor d(852) xor d(850) xor d(849) xor d(846) xor d(838) xor d(837) xor d(836) xor d(835) xor d(831) xor d(830) xor d(829) xor d(827) xor d(826) xor d(823) xor d(821) xor d(820) xor d(819) xor d(818) xor d(816) xor d(815) xor d(808) xor d(807) xor d(805) xor d(804) xor d(803) xor d(801) xor d(799) xor d(798) xor d(797) xor d(796) xor d(795) xor d(790) xor d(788) xor d(787) xor d(784) xor d(782) xor d(780) xor d(779) xor d(778) xor d(774) xor d(772) xor d(771) xor d(770) xor d(769) xor d(766) xor d(765) xor d(761) xor d(757) xor d(754) xor d(752) xor d(751) xor d(749) xor d(745) xor d(744) xor d(743) xor d(742) xor d(741) xor d(738) xor d(737) xor d(735) xor d(733) xor d(729) xor d(728) xor d(727) xor d(724) xor d(723) xor d(722) xor d(720) xor d(718) xor d(717) xor d(716) xor d(715) xor d(713) xor d(712) xor d(711) xor d(710) xor d(705) xor d(704) xor d(702) xor d(700) xor d(697) xor d(696) xor d(695) xor d(694) xor d(692) xor d(691) xor d(690) xor d(688) xor d(686) xor d(683) xor d(682) xor d(681) xor d(680) xor d(676) xor d(675) xor d(674) xor d(672) xor d(669) xor d(668) xor d(667) xor d(666) xor d(664) xor d(663) xor d(662) xor d(661) xor d(660) xor d(659) xor d(658) xor d(656) xor d(652) xor d(650) xor d(648) xor d(644) xor d(643) xor d(640) xor d(638) xor d(637) xor d(636) xor d(635) xor d(631) xor d(628) xor d(624) xor d(621) xor d(620) xor d(619) xor d(615) xor d(614) xor d(613) xor d(612) xor d(611) xor d(610) xor d(609) xor d(605) xor d(602) xor d(601) xor d(599) xor d(598) xor d(597) xor d(594) xor d(592) xor d(591) xor d(590) xor d(589) xor d(588) xor d(586) xor d(585) xor d(583) xor d(582) xor d(579) xor d(578) xor d(575) xor d(573) xor d(572) xor d(571) xor d(569) xor d(568) xor d(567) xor d(564) xor d(562) xor d(561) xor d(560) xor d(558) xor d(557) xor d(554) xor d(550) xor d(548) xor d(547) xor d(546) xor d(544) xor d(543) xor d(542) xor d(540) xor d(539) xor d(538) xor d(532) xor d(529) xor d(528) xor d(527) xor d(524) xor d(523) xor d(522) xor d(519) xor d(517) xor d(515) xor d(510) xor d(508) xor d(507) xor d(506) xor d(505) xor d(504) xor d(501) xor d(500) xor d(496) xor d(495) xor d(493) xor d(492) xor d(488) xor d(487) xor d(486) xor d(484) xor d(477) xor d(476) xor d(473) xor d(472) xor d(471) xor d(470) xor d(466) xor d(464) xor d(462) xor d(461) xor d(460) xor d(458) xor d(457) xor d(455) xor d(453) xor d(451) xor d(450) xor d(446) xor d(444) xor d(437) xor d(436) xor d(435) xor d(430) xor d(428) xor d(427) xor d(425) xor d(423) xor d(419) xor d(418) xor d(417) xor d(416) xor d(415) xor d(414) xor d(411) xor d(409) xor d(407) xor d(406) xor d(405) xor d(402) xor d(396) xor d(395) xor d(394) xor d(391) xor d(387) xor d(386) xor d(385) xor d(384) xor d(380) xor d(379) xor d(378) xor d(375) xor d(372) xor d(370) xor d(368) xor d(367) xor d(364) xor d(363) xor d(362) xor d(360) xor d(358) xor d(357) xor d(355) xor d(354) xor d(351) xor d(341) xor d(340) xor d(339) xor d(336) xor d(335) xor d(332) xor d(330) xor d(329) xor d(326) xor d(325) xor d(324) xor d(320) xor d(318) xor d(314) xor d(313) xor d(312) xor d(311) xor d(308) xor d(306) xor d(305) xor d(303) xor d(297) xor d(291) xor d(290) xor d(280) xor d(279) xor d(278) xor d(277) xor d(275) xor d(273) xor d(269) xor d(266) xor d(265) xor d(261) xor d(259) xor d(257) xor d(256) xor d(255) xor d(253) xor d(251) xor d(248) xor d(246) xor d(245) xor d(244) xor d(243) xor d(242) xor d(241) xor d(235) xor d(234) xor d(230) xor d(229) xor d(228) xor d(227) xor d(222) xor d(220) xor d(219) xor d(218) xor d(217) xor d(216) xor d(215) xor d(214) xor d(210) xor d(207) xor d(206) xor d(204) xor d(201) xor d(199) xor d(197) xor d(196) xor d(194) xor d(193) xor d(192) xor d(190) xor d(188) xor d(187) xor d(185) xor d(184) xor d(181) xor d(180) xor d(177) xor d(175) xor d(170) xor d(169) xor d(168) xor d(167) xor d(165) xor d(162) xor d(158) xor d(157) xor d(156) xor d(154) xor d(153) xor d(149) xor d(145) xor d(141) xor d(137) xor d(136) xor d(134) xor d(133) xor d(128) xor d(127) xor d(122) xor d(121) xor d(120) xor d(119) xor d(117) xor d(116) xor d(113) xor d(111) xor d(110) xor d(109) xor d(108) xor d(105) xor d(102) xor d(101) xor d(98) xor d(97) xor d(96) xor d(94) xor d(92) xor d(91) xor d(87) xor d(86) xor d(85) xor d(82) xor d(81) xor d(77) xor d(75) xor d(74) xor d(73) xor d(71) xor d(69) xor d(68) xor d(63) xor d(61) xor d(59) xor d(57) xor d(56) xor d(54) xor d(53) xor d(52) xor d(51) xor d(50) xor d(49) xor d(47) xor d(46) xor d(42) xor d(41) xor d(31) xor d(30) xor d(27) xor d(24) xor d(21) xor d(18) xor d(17) xor d(15) xor d(13) xor d(12) xor d(9) xor d(6) xor d(5) xor d(4) xor d(2) xor d(1) xor d(0) xor c(0) xor c(1) xor c(3) xor c(4) xor c(9) xor c(10) xor c(13) xor c(14) xor c(15) xor c(18) xor c(23) xor c(24) xor c(26) xor c(27) xor c(28) xor c(29) xor c(30) xor c(31);
    newcrc(13) := d(1023) xor d(1022) xor d(1021) xor d(1020) xor d(1019) xor d(1017) xor d(1016) xor d(1011) xor d(1008) xor d(1007) xor d(1006) xor d(1003) xor d(1002) xor d(997) xor d(996) xor d(994) xor d(993) xor d(991) xor d(990) xor d(988) xor d(986) xor d(985) xor d(984) xor d(980) xor d(979) xor d(978) xor d(977) xor d(974) xor d(973) xor d(971) xor d(970) xor d(969) xor d(966) xor d(963) xor d(962) xor d(961) xor d(960) xor d(959) xor d(958) xor d(954) xor d(950) xor d(943) xor d(942) xor d(940) xor d(937) xor d(929) xor d(928) xor d(923) xor d(922) xor d(919) xor d(918) xor d(917) xor d(916) xor d(911) xor d(910) xor d(909) xor d(907) xor d(906) xor d(903) xor d(902) xor d(901) xor d(898) xor d(896) xor d(889) xor d(888) xor d(887) xor d(886) xor d(881) xor d(880) xor d(876) xor d(875) xor d(873) xor d(872) xor d(871) xor d(868) xor d(867) xor d(864) xor d(862) xor d(859) xor d(858) xor d(857) xor d(856) xor d(853) xor d(851) xor d(850) xor d(847) xor d(839) xor d(838) xor d(837) xor d(836) xor d(832) xor d(831) xor d(830) xor d(828) xor d(827) xor d(824) xor d(822) xor d(821) xor d(820) xor d(819) xor d(817) xor d(816) xor d(809) xor d(808) xor d(806) xor d(805) xor d(804) xor d(802) xor d(800) xor d(799) xor d(798) xor d(797) xor d(796) xor d(791) xor d(789) xor d(788) xor d(785) xor d(783) xor d(781) xor d(780) xor d(779) xor d(775) xor d(773) xor d(772) xor d(771) xor d(770) xor d(767) xor d(766) xor d(762) xor d(758) xor d(755) xor d(753) xor d(752) xor d(750) xor d(746) xor d(745) xor d(744) xor d(743) xor d(742) xor d(739) xor d(738) xor d(736) xor d(734) xor d(730) xor d(729) xor d(728) xor d(725) xor d(724) xor d(723) xor d(721) xor d(719) xor d(718) xor d(717) xor d(716) xor d(714) xor d(713) xor d(712) xor d(711) xor d(706) xor d(705) xor d(703) xor d(701) xor d(698) xor d(697) xor d(696) xor d(695) xor d(693) xor d(692) xor d(691) xor d(689) xor d(687) xor d(684) xor d(683) xor d(682) xor d(681) xor d(677) xor d(676) xor d(675) xor d(673) xor d(670) xor d(669) xor d(668) xor d(667) xor d(665) xor d(664) xor d(663) xor d(662) xor d(661) xor d(660) xor d(659) xor d(657) xor d(653) xor d(651) xor d(649) xor d(645) xor d(644) xor d(641) xor d(639) xor d(638) xor d(637) xor d(636) xor d(632) xor d(629) xor d(625) xor d(622) xor d(621) xor d(620) xor d(616) xor d(615) xor d(614) xor d(613) xor d(612) xor d(611) xor d(610) xor d(606) xor d(603) xor d(602) xor d(600) xor d(599) xor d(598) xor d(595) xor d(593) xor d(592) xor d(591) xor d(590) xor d(589) xor d(587) xor d(586) xor d(584) xor d(583) xor d(580) xor d(579) xor d(576) xor d(574) xor d(573) xor d(572) xor d(570) xor d(569) xor d(568) xor d(565) xor d(563) xor d(562) xor d(561) xor d(559) xor d(558) xor d(555) xor d(551) xor d(549) xor d(548) xor d(547) xor d(545) xor d(544) xor d(543) xor d(541) xor d(540) xor d(539) xor d(533) xor d(530) xor d(529) xor d(528) xor d(525) xor d(524) xor d(523) xor d(520) xor d(518) xor d(516) xor d(511) xor d(509) xor d(508) xor d(507) xor d(506) xor d(505) xor d(502) xor d(501) xor d(497) xor d(496) xor d(494) xor d(493) xor d(489) xor d(488) xor d(487) xor d(485) xor d(478) xor d(477) xor d(474) xor d(473) xor d(472) xor d(471) xor d(467) xor d(465) xor d(463) xor d(462) xor d(461) xor d(459) xor d(458) xor d(456) xor d(454) xor d(452) xor d(451) xor d(447) xor d(445) xor d(438) xor d(437) xor d(436) xor d(431) xor d(429) xor d(428) xor d(426) xor d(424) xor d(420) xor d(419) xor d(418) xor d(417) xor d(416) xor d(415) xor d(412) xor d(410) xor d(408) xor d(407) xor d(406) xor d(403) xor d(397) xor d(396) xor d(395) xor d(392) xor d(388) xor d(387) xor d(386) xor d(385) xor d(381) xor d(380) xor d(379) xor d(376) xor d(373) xor d(371) xor d(369) xor d(368) xor d(365) xor d(364) xor d(363) xor d(361) xor d(359) xor d(358) xor d(356) xor d(355) xor d(352) xor d(342) xor d(341) xor d(340) xor d(337) xor d(336) xor d(333) xor d(331) xor d(330) xor d(327) xor d(326) xor d(325) xor d(321) xor d(319) xor d(315) xor d(314) xor d(313) xor d(312) xor d(309) xor d(307) xor d(306) xor d(304) xor d(298) xor d(292) xor d(291) xor d(281) xor d(280) xor d(279) xor d(278) xor d(276) xor d(274) xor d(270) xor d(267) xor d(266) xor d(262) xor d(260) xor d(258) xor d(257) xor d(256) xor d(254) xor d(252) xor d(249) xor d(247) xor d(246) xor d(245) xor d(244) xor d(243) xor d(242) xor d(236) xor d(235) xor d(231) xor d(230) xor d(229) xor d(228) xor d(223) xor d(221) xor d(220) xor d(219) xor d(218) xor d(217) xor d(216) xor d(215) xor d(211) xor d(208) xor d(207) xor d(205) xor d(202) xor d(200) xor d(198) xor d(197) xor d(195) xor d(194) xor d(193) xor d(191) xor d(189) xor d(188) xor d(186) xor d(185) xor d(182) xor d(181) xor d(178) xor d(176) xor d(171) xor d(170) xor d(169) xor d(168) xor d(166) xor d(163) xor d(159) xor d(158) xor d(157) xor d(155) xor d(154) xor d(150) xor d(146) xor d(142) xor d(138) xor d(137) xor d(135) xor d(134) xor d(129) xor d(128) xor d(123) xor d(122) xor d(121) xor d(120) xor d(118) xor d(117) xor d(114) xor d(112) xor d(111) xor d(110) xor d(109) xor d(106) xor d(103) xor d(102) xor d(99) xor d(98) xor d(97) xor d(95) xor d(93) xor d(92) xor d(88) xor d(87) xor d(86) xor d(83) xor d(82) xor d(78) xor d(76) xor d(75) xor d(74) xor d(72) xor d(70) xor d(69) xor d(64) xor d(62) xor d(60) xor d(58) xor d(57) xor d(55) xor d(54) xor d(53) xor d(52) xor d(51) xor d(50) xor d(48) xor d(47) xor d(43) xor d(42) xor d(32) xor d(31) xor d(28) xor d(25) xor d(22) xor d(19) xor d(18) xor d(16) xor d(14) xor d(13) xor d(10) xor d(7) xor d(6) xor d(5) xor d(3) xor d(2) xor d(1) xor c(1) xor c(2) xor c(4) xor c(5) xor c(10) xor c(11) xor c(14) xor c(15) xor c(16) xor c(19) xor c(24) xor c(25) xor c(27) xor c(28) xor c(29) xor c(30) xor c(31);
    newcrc(14) := d(1023) xor d(1022) xor d(1021) xor d(1020) xor d(1018) xor d(1017) xor d(1012) xor d(1009) xor d(1008) xor d(1007) xor d(1004) xor d(1003) xor d(998) xor d(997) xor d(995) xor d(994) xor d(992) xor d(991) xor d(989) xor d(987) xor d(986) xor d(985) xor d(981) xor d(980) xor d(979) xor d(978) xor d(975) xor d(974) xor d(972) xor d(971) xor d(970) xor d(967) xor d(964) xor d(963) xor d(962) xor d(961) xor d(960) xor d(959) xor d(955) xor d(951) xor d(944) xor d(943) xor d(941) xor d(938) xor d(930) xor d(929) xor d(924) xor d(923) xor d(920) xor d(919) xor d(918) xor d(917) xor d(912) xor d(911) xor d(910) xor d(908) xor d(907) xor d(904) xor d(903) xor d(902) xor d(899) xor d(897) xor d(890) xor d(889) xor d(888) xor d(887) xor d(882) xor d(881) xor d(877) xor d(876) xor d(874) xor d(873) xor d(872) xor d(869) xor d(868) xor d(865) xor d(863) xor d(860) xor d(859) xor d(858) xor d(857) xor d(854) xor d(852) xor d(851) xor d(848) xor d(840) xor d(839) xor d(838) xor d(837) xor d(833) xor d(832) xor d(831) xor d(829) xor d(828) xor d(825) xor d(823) xor d(822) xor d(821) xor d(820) xor d(818) xor d(817) xor d(810) xor d(809) xor d(807) xor d(806) xor d(805) xor d(803) xor d(801) xor d(800) xor d(799) xor d(798) xor d(797) xor d(792) xor d(790) xor d(789) xor d(786) xor d(784) xor d(782) xor d(781) xor d(780) xor d(776) xor d(774) xor d(773) xor d(772) xor d(771) xor d(768) xor d(767) xor d(763) xor d(759) xor d(756) xor d(754) xor d(753) xor d(751) xor d(747) xor d(746) xor d(745) xor d(744) xor d(743) xor d(740) xor d(739) xor d(737) xor d(735) xor d(731) xor d(730) xor d(729) xor d(726) xor d(725) xor d(724) xor d(722) xor d(720) xor d(719) xor d(718) xor d(717) xor d(715) xor d(714) xor d(713) xor d(712) xor d(707) xor d(706) xor d(704) xor d(702) xor d(699) xor d(698) xor d(697) xor d(696) xor d(694) xor d(693) xor d(692) xor d(690) xor d(688) xor d(685) xor d(684) xor d(683) xor d(682) xor d(678) xor d(677) xor d(676) xor d(674) xor d(671) xor d(670) xor d(669) xor d(668) xor d(666) xor d(665) xor d(664) xor d(663) xor d(662) xor d(661) xor d(660) xor d(658) xor d(654) xor d(652) xor d(650) xor d(646) xor d(645) xor d(642) xor d(640) xor d(639) xor d(638) xor d(637) xor d(633) xor d(630) xor d(626) xor d(623) xor d(622) xor d(621) xor d(617) xor d(616) xor d(615) xor d(614) xor d(613) xor d(612) xor d(611) xor d(607) xor d(604) xor d(603) xor d(601) xor d(600) xor d(599) xor d(596) xor d(594) xor d(593) xor d(592) xor d(591) xor d(590) xor d(588) xor d(587) xor d(585) xor d(584) xor d(581) xor d(580) xor d(577) xor d(575) xor d(574) xor d(573) xor d(571) xor d(570) xor d(569) xor d(566) xor d(564) xor d(563) xor d(562) xor d(560) xor d(559) xor d(556) xor d(552) xor d(550) xor d(549) xor d(548) xor d(546) xor d(545) xor d(544) xor d(542) xor d(541) xor d(540) xor d(534) xor d(531) xor d(530) xor d(529) xor d(526) xor d(525) xor d(524) xor d(521) xor d(519) xor d(517) xor d(512) xor d(510) xor d(509) xor d(508) xor d(507) xor d(506) xor d(503) xor d(502) xor d(498) xor d(497) xor d(495) xor d(494) xor d(490) xor d(489) xor d(488) xor d(486) xor d(479) xor d(478) xor d(475) xor d(474) xor d(473) xor d(472) xor d(468) xor d(466) xor d(464) xor d(463) xor d(462) xor d(460) xor d(459) xor d(457) xor d(455) xor d(453) xor d(452) xor d(448) xor d(446) xor d(439) xor d(438) xor d(437) xor d(432) xor d(430) xor d(429) xor d(427) xor d(425) xor d(421) xor d(420) xor d(419) xor d(418) xor d(417) xor d(416) xor d(413) xor d(411) xor d(409) xor d(408) xor d(407) xor d(404) xor d(398) xor d(397) xor d(396) xor d(393) xor d(389) xor d(388) xor d(387) xor d(386) xor d(382) xor d(381) xor d(380) xor d(377) xor d(374) xor d(372) xor d(370) xor d(369) xor d(366) xor d(365) xor d(364) xor d(362) xor d(360) xor d(359) xor d(357) xor d(356) xor d(353) xor d(343) xor d(342) xor d(341) xor d(338) xor d(337) xor d(334) xor d(332) xor d(331) xor d(328) xor d(327) xor d(326) xor d(322) xor d(320) xor d(316) xor d(315) xor d(314) xor d(313) xor d(310) xor d(308) xor d(307) xor d(305) xor d(299) xor d(293) xor d(292) xor d(282) xor d(281) xor d(280) xor d(279) xor d(277) xor d(275) xor d(271) xor d(268) xor d(267) xor d(263) xor d(261) xor d(259) xor d(258) xor d(257) xor d(255) xor d(253) xor d(250) xor d(248) xor d(247) xor d(246) xor d(245) xor d(244) xor d(243) xor d(237) xor d(236) xor d(232) xor d(231) xor d(230) xor d(229) xor d(224) xor d(222) xor d(221) xor d(220) xor d(219) xor d(218) xor d(217) xor d(216) xor d(212) xor d(209) xor d(208) xor d(206) xor d(203) xor d(201) xor d(199) xor d(198) xor d(196) xor d(195) xor d(194) xor d(192) xor d(190) xor d(189) xor d(187) xor d(186) xor d(183) xor d(182) xor d(179) xor d(177) xor d(172) xor d(171) xor d(170) xor d(169) xor d(167) xor d(164) xor d(160) xor d(159) xor d(158) xor d(156) xor d(155) xor d(151) xor d(147) xor d(143) xor d(139) xor d(138) xor d(136) xor d(135) xor d(130) xor d(129) xor d(124) xor d(123) xor d(122) xor d(121) xor d(119) xor d(118) xor d(115) xor d(113) xor d(112) xor d(111) xor d(110) xor d(107) xor d(104) xor d(103) xor d(100) xor d(99) xor d(98) xor d(96) xor d(94) xor d(93) xor d(89) xor d(88) xor d(87) xor d(84) xor d(83) xor d(79) xor d(77) xor d(76) xor d(75) xor d(73) xor d(71) xor d(70) xor d(65) xor d(63) xor d(61) xor d(59) xor d(58) xor d(56) xor d(55) xor d(54) xor d(53) xor d(52) xor d(51) xor d(49) xor d(48) xor d(44) xor d(43) xor d(33) xor d(32) xor d(29) xor d(26) xor d(23) xor d(20) xor d(19) xor d(17) xor d(15) xor d(14) xor d(11) xor d(8) xor d(7) xor d(6) xor d(4) xor d(3) xor d(2) xor c(0) xor c(2) xor c(3) xor c(5) xor c(6) xor c(11) xor c(12) xor c(15) xor c(16) xor c(17) xor c(20) xor c(25) xor c(26) xor c(28) xor c(29) xor c(30) xor c(31);
    newcrc(15) := d(1023) xor d(1022) xor d(1021) xor d(1019) xor d(1018) xor d(1013) xor d(1010) xor d(1009) xor d(1008) xor d(1005) xor d(1004) xor d(999) xor d(998) xor d(996) xor d(995) xor d(993) xor d(992) xor d(990) xor d(988) xor d(987) xor d(986) xor d(982) xor d(981) xor d(980) xor d(979) xor d(976) xor d(975) xor d(973) xor d(972) xor d(971) xor d(968) xor d(965) xor d(964) xor d(963) xor d(962) xor d(961) xor d(960) xor d(956) xor d(952) xor d(945) xor d(944) xor d(942) xor d(939) xor d(931) xor d(930) xor d(925) xor d(924) xor d(921) xor d(920) xor d(919) xor d(918) xor d(913) xor d(912) xor d(911) xor d(909) xor d(908) xor d(905) xor d(904) xor d(903) xor d(900) xor d(898) xor d(891) xor d(890) xor d(889) xor d(888) xor d(883) xor d(882) xor d(878) xor d(877) xor d(875) xor d(874) xor d(873) xor d(870) xor d(869) xor d(866) xor d(864) xor d(861) xor d(860) xor d(859) xor d(858) xor d(855) xor d(853) xor d(852) xor d(849) xor d(841) xor d(840) xor d(839) xor d(838) xor d(834) xor d(833) xor d(832) xor d(830) xor d(829) xor d(826) xor d(824) xor d(823) xor d(822) xor d(821) xor d(819) xor d(818) xor d(811) xor d(810) xor d(808) xor d(807) xor d(806) xor d(804) xor d(802) xor d(801) xor d(800) xor d(799) xor d(798) xor d(793) xor d(791) xor d(790) xor d(787) xor d(785) xor d(783) xor d(782) xor d(781) xor d(777) xor d(775) xor d(774) xor d(773) xor d(772) xor d(769) xor d(768) xor d(764) xor d(760) xor d(757) xor d(755) xor d(754) xor d(752) xor d(748) xor d(747) xor d(746) xor d(745) xor d(744) xor d(741) xor d(740) xor d(738) xor d(736) xor d(732) xor d(731) xor d(730) xor d(727) xor d(726) xor d(725) xor d(723) xor d(721) xor d(720) xor d(719) xor d(718) xor d(716) xor d(715) xor d(714) xor d(713) xor d(708) xor d(707) xor d(705) xor d(703) xor d(700) xor d(699) xor d(698) xor d(697) xor d(695) xor d(694) xor d(693) xor d(691) xor d(689) xor d(686) xor d(685) xor d(684) xor d(683) xor d(679) xor d(678) xor d(677) xor d(675) xor d(672) xor d(671) xor d(670) xor d(669) xor d(667) xor d(666) xor d(665) xor d(664) xor d(663) xor d(662) xor d(661) xor d(659) xor d(655) xor d(653) xor d(651) xor d(647) xor d(646) xor d(643) xor d(641) xor d(640) xor d(639) xor d(638) xor d(634) xor d(631) xor d(627) xor d(624) xor d(623) xor d(622) xor d(618) xor d(617) xor d(616) xor d(615) xor d(614) xor d(613) xor d(612) xor d(608) xor d(605) xor d(604) xor d(602) xor d(601) xor d(600) xor d(597) xor d(595) xor d(594) xor d(593) xor d(592) xor d(591) xor d(589) xor d(588) xor d(586) xor d(585) xor d(582) xor d(581) xor d(578) xor d(576) xor d(575) xor d(574) xor d(572) xor d(571) xor d(570) xor d(567) xor d(565) xor d(564) xor d(563) xor d(561) xor d(560) xor d(557) xor d(553) xor d(551) xor d(550) xor d(549) xor d(547) xor d(546) xor d(545) xor d(543) xor d(542) xor d(541) xor d(535) xor d(532) xor d(531) xor d(530) xor d(527) xor d(526) xor d(525) xor d(522) xor d(520) xor d(518) xor d(513) xor d(511) xor d(510) xor d(509) xor d(508) xor d(507) xor d(504) xor d(503) xor d(499) xor d(498) xor d(496) xor d(495) xor d(491) xor d(490) xor d(489) xor d(487) xor d(480) xor d(479) xor d(476) xor d(475) xor d(474) xor d(473) xor d(469) xor d(467) xor d(465) xor d(464) xor d(463) xor d(461) xor d(460) xor d(458) xor d(456) xor d(454) xor d(453) xor d(449) xor d(447) xor d(440) xor d(439) xor d(438) xor d(433) xor d(431) xor d(430) xor d(428) xor d(426) xor d(422) xor d(421) xor d(420) xor d(419) xor d(418) xor d(417) xor d(414) xor d(412) xor d(410) xor d(409) xor d(408) xor d(405) xor d(399) xor d(398) xor d(397) xor d(394) xor d(390) xor d(389) xor d(388) xor d(387) xor d(383) xor d(382) xor d(381) xor d(378) xor d(375) xor d(373) xor d(371) xor d(370) xor d(367) xor d(366) xor d(365) xor d(363) xor d(361) xor d(360) xor d(358) xor d(357) xor d(354) xor d(344) xor d(343) xor d(342) xor d(339) xor d(338) xor d(335) xor d(333) xor d(332) xor d(329) xor d(328) xor d(327) xor d(323) xor d(321) xor d(317) xor d(316) xor d(315) xor d(314) xor d(311) xor d(309) xor d(308) xor d(306) xor d(300) xor d(294) xor d(293) xor d(283) xor d(282) xor d(281) xor d(280) xor d(278) xor d(276) xor d(272) xor d(269) xor d(268) xor d(264) xor d(262) xor d(260) xor d(259) xor d(258) xor d(256) xor d(254) xor d(251) xor d(249) xor d(248) xor d(247) xor d(246) xor d(245) xor d(244) xor d(238) xor d(237) xor d(233) xor d(232) xor d(231) xor d(230) xor d(225) xor d(223) xor d(222) xor d(221) xor d(220) xor d(219) xor d(218) xor d(217) xor d(213) xor d(210) xor d(209) xor d(207) xor d(204) xor d(202) xor d(200) xor d(199) xor d(197) xor d(196) xor d(195) xor d(193) xor d(191) xor d(190) xor d(188) xor d(187) xor d(184) xor d(183) xor d(180) xor d(178) xor d(173) xor d(172) xor d(171) xor d(170) xor d(168) xor d(165) xor d(161) xor d(160) xor d(159) xor d(157) xor d(156) xor d(152) xor d(148) xor d(144) xor d(140) xor d(139) xor d(137) xor d(136) xor d(131) xor d(130) xor d(125) xor d(124) xor d(123) xor d(122) xor d(120) xor d(119) xor d(116) xor d(114) xor d(113) xor d(112) xor d(111) xor d(108) xor d(105) xor d(104) xor d(101) xor d(100) xor d(99) xor d(97) xor d(95) xor d(94) xor d(90) xor d(89) xor d(88) xor d(85) xor d(84) xor d(80) xor d(78) xor d(77) xor d(76) xor d(74) xor d(72) xor d(71) xor d(66) xor d(64) xor d(62) xor d(60) xor d(59) xor d(57) xor d(56) xor d(55) xor d(54) xor d(53) xor d(52) xor d(50) xor d(49) xor d(45) xor d(44) xor d(34) xor d(33) xor d(30) xor d(27) xor d(24) xor d(21) xor d(20) xor d(18) xor d(16) xor d(15) xor d(12) xor d(9) xor d(8) xor d(7) xor d(5) xor d(4) xor d(3) xor c(0) xor c(1) xor c(3) xor c(4) xor c(6) xor c(7) xor c(12) xor c(13) xor c(16) xor c(17) xor c(18) xor c(21) xor c(26) xor c(27) xor c(29) xor c(30) xor c(31);
    newcrc(16) := d(1023) xor d(1022) xor d(1021) xor d(1020) xor d(1018) xor d(1016) xor d(1015) xor d(1014) xor d(1012) xor d(1010) xor d(1008) xor d(1004) xor d(998) xor d(997) xor d(993) xor d(992) xor d(991) xor d(990) xor d(989) xor d(988) xor d(987) xor d(985) xor d(984) xor d(979) xor d(978) xor d(976) xor d(975) xor d(973) xor d(972) xor d(971) xor d(969) xor d(967) xor d(966) xor d(965) xor d(964) xor d(963) xor d(962) xor d(961) xor d(960) xor d(959) xor d(958) xor d(957) xor d(955) xor d(954) xor d(950) xor d(948) xor d(946) xor d(945) xor d(944) xor d(943) xor d(941) xor d(940) xor d(939) xor d(938) xor d(935) xor d(934) xor d(933) xor d(932) xor d(926) xor d(925) xor d(922) xor d(921) xor d(919) xor d(918) xor d(917) xor d(915) xor d(914) xor d(913) xor d(912) xor d(909) xor d(907) xor d(905) xor d(903) xor d(902) xor d(900) xor d(898) xor d(897) xor d(896) xor d(893) xor d(892) xor d(887) xor d(886) xor d(884) xor d(881) xor d(877) xor d(873) xor d(870) xor d(869) xor d(868) xor d(865) xor d(863) xor d(862) xor d(857) xor d(856) xor d(851) xor d(849) xor d(848) xor d(846) xor d(841) xor d(837) xor d(833) xor d(832) xor d(831) xor d(830) xor d(823) xor d(822) xor d(820) xor d(818) xor d(816) xor d(815) xor d(814) xor d(813) xor d(810) xor d(806) xor d(805) xor d(804) xor d(801) xor d(799) xor d(798) xor d(794) xor d(793) xor d(792) xor d(785) xor d(783) xor d(780) xor d(778) xor d(775) xor d(773) xor d(770) xor d(767) xor d(763) xor d(762) xor d(761) xor d(750) xor d(749) xor d(746) xor d(745) xor d(744) xor d(740) xor d(739) xor d(737) xor d(736) xor d(733) xor d(729) xor d(728) xor d(726) xor d(725) xor d(723) xor d(717) xor d(716) xor d(714) xor d(710) xor d(709) xor d(707) xor d(706) xor d(702) xor d(699) xor d(696) xor d(693) xor d(692) xor d(691) xor d(690) xor d(689) xor d(685) xor d(684) xor d(679) xor d(678) xor d(676) xor d(675) xor d(674) xor d(671) xor d(669) xor d(664) xor d(663) xor d(662) xor d(660) xor d(658) xor d(655) xor d(654) xor d(653) xor d(649) xor d(647) xor d(646) xor d(641) xor d(639) xor d(636) xor d(635) xor d(630) xor d(629) xor d(628) xor d(626) xor d(625) xor d(620) xor d(618) xor d(616) xor d(614) xor d(612) xor d(611) xor d(610) xor d(607) xor d(605) xor d(604) xor d(601) xor d(600) xor d(599) xor d(598) xor d(594) xor d(591) xor d(590) xor d(589) xor d(585) xor d(582) xor d(580) xor d(579) xor d(578) xor d(577) xor d(576) xor d(574) xor d(572) xor d(568) xor d(567) xor d(566) xor d(564) xor d(563) xor d(562) xor d(560) xor d(557) xor d(556) xor d(555) xor d(552) xor d(550) xor d(549) xor d(548) xor d(547) xor d(546) xor d(545) xor d(544) xor d(543) xor d(540) xor d(539) xor d(536) xor d(535) xor d(534) xor d(533) xor d(530) xor d(529) xor d(527) xor d(525) xor d(523) xor d(522) xor d(518) xor d(516) xor d(509) xor d(507) xor d(506) xor d(505) xor d(504) xor d(502) xor d(501) xor d(499) xor d(497) xor d(496) xor d(495) xor d(494) xor d(493) xor d(489) xor d(486) xor d(483) xor d(482) xor d(479) xor d(475) xor d(474) xor d(472) xor d(466) xor d(459) xor d(458) xor d(457) xor d(455) xor d(454) xor d(452) xor d(449) xor d(444) xor d(441) xor d(440) xor d(439) xor d(437) xor d(436) xor d(433) xor d(432) xor d(431) xor d(429) xor d(427) xor d(424) xor d(423) xor d(421) xor d(420) xor d(416) xor d(415) xor d(414) xor d(413) xor d(412) xor d(411) xor d(410) xor d(408) xor d(407) xor d(406) xor d(405) xor d(404) xor d(396) xor d(395) xor d(393) xor d(392) xor d(389) xor d(387) xor d(386) xor d(384) xor d(383) xor d(382) xor d(381) xor d(379) xor d(378) xor d(371) xor d(369) xor d(367) xor d(364) xor d(363) xor d(361) xor d(357) xor d(355) xor d(353) xor d(349) xor d(348) xor d(347) xor d(343) xor d(342) xor d(341) xor d(340) xor d(338) xor d(337) xor d(336) xor d(335) xor d(330) xor d(329) xor d(327) xor d(324) xor d(321) xor d(320) xor d(319) xor d(316) xor d(307) xor d(305) xor d(303) xor d(302) xor d(301) xor d(300) xor d(299) xor d(298) xor d(297) xor d(296) xor d(292) xor d(290) xor d(288) xor d(287) xor d(286) xor d(284) xor d(282) xor d(281) xor d(276) xor d(274) xor d(270) xor d(268) xor d(264) xor d(263) xor d(260) xor d(250) xor d(249) xor d(247) xor d(246) xor d(245) xor d(243) xor d(239) xor d(238) xor d(237) xor d(233) xor d(232) xor d(231) xor d(230) xor d(228) xor d(227) xor d(223) xor d(222) xor d(221) xor d(220) xor d(219) xor d(218) xor d(216) xor d(212) xor d(211) xor d(209) xor d(207) xor d(205) xor d(202) xor d(200) xor d(199) xor d(196) xor d(193) xor d(190) xor d(189) xor d(186) xor d(185) xor d(184) xor d(183) xor d(182) xor d(181) xor d(179) xor d(174) xor d(173) xor d(170) xor d(167) xor d(160) xor d(157) xor d(156) xor d(155) xor d(153) xor d(151) xor d(145) xor d(144) xor d(143) xor d(141) xor d(140) xor d(138) xor d(136) xor d(135) xor d(134) xor d(131) xor d(128) xor d(127) xor d(124) xor d(121) xor d(120) xor d(119) xor d(118) xor d(116) xor d(115) xor d(112) xor d(111) xor d(110) xor d(109) xor d(105) xor d(104) xor d(103) xor d(102) xor d(100) xor d(99) xor d(97) xor d(94) xor d(91) xor d(90) xor d(89) xor d(87) xor d(86) xor d(84) xor d(83) xor d(82) xor d(78) xor d(77) xor d(75) xor d(68) xor d(66) xor d(57) xor d(56) xor d(51) xor d(48) xor d(47) xor d(46) xor d(44) xor d(37) xor d(35) xor d(32) xor d(30) xor d(29) xor d(26) xor d(24) xor d(22) xor d(21) xor d(19) xor d(17) xor d(13) xor d(12) xor d(8) xor d(5) xor d(4) xor d(0) xor c(0) xor c(1) xor c(5) xor c(6) xor c(12) xor c(16) xor c(18) xor c(20) xor c(22) xor c(23) xor c(24) xor c(26) xor c(28) xor c(29) xor c(30) xor c(31);
    newcrc(17) := d(1023) xor d(1022) xor d(1021) xor d(1019) xor d(1017) xor d(1016) xor d(1015) xor d(1013) xor d(1011) xor d(1009) xor d(1005) xor d(999) xor d(998) xor d(994) xor d(993) xor d(992) xor d(991) xor d(990) xor d(989) xor d(988) xor d(986) xor d(985) xor d(980) xor d(979) xor d(977) xor d(976) xor d(974) xor d(973) xor d(972) xor d(970) xor d(968) xor d(967) xor d(966) xor d(965) xor d(964) xor d(963) xor d(962) xor d(961) xor d(960) xor d(959) xor d(958) xor d(956) xor d(955) xor d(951) xor d(949) xor d(947) xor d(946) xor d(945) xor d(944) xor d(942) xor d(941) xor d(940) xor d(939) xor d(936) xor d(935) xor d(934) xor d(933) xor d(927) xor d(926) xor d(923) xor d(922) xor d(920) xor d(919) xor d(918) xor d(916) xor d(915) xor d(914) xor d(913) xor d(910) xor d(908) xor d(906) xor d(904) xor d(903) xor d(901) xor d(899) xor d(898) xor d(897) xor d(894) xor d(893) xor d(888) xor d(887) xor d(885) xor d(882) xor d(878) xor d(874) xor d(871) xor d(870) xor d(869) xor d(866) xor d(864) xor d(863) xor d(858) xor d(857) xor d(852) xor d(850) xor d(849) xor d(847) xor d(842) xor d(838) xor d(834) xor d(833) xor d(832) xor d(831) xor d(824) xor d(823) xor d(821) xor d(819) xor d(817) xor d(816) xor d(815) xor d(814) xor d(811) xor d(807) xor d(806) xor d(805) xor d(802) xor d(800) xor d(799) xor d(795) xor d(794) xor d(793) xor d(786) xor d(784) xor d(781) xor d(779) xor d(776) xor d(774) xor d(771) xor d(768) xor d(764) xor d(763) xor d(762) xor d(751) xor d(750) xor d(747) xor d(746) xor d(745) xor d(741) xor d(740) xor d(738) xor d(737) xor d(734) xor d(730) xor d(729) xor d(727) xor d(726) xor d(724) xor d(718) xor d(717) xor d(715) xor d(711) xor d(710) xor d(708) xor d(707) xor d(703) xor d(700) xor d(697) xor d(694) xor d(693) xor d(692) xor d(691) xor d(690) xor d(686) xor d(685) xor d(680) xor d(679) xor d(677) xor d(676) xor d(675) xor d(672) xor d(670) xor d(665) xor d(664) xor d(663) xor d(661) xor d(659) xor d(656) xor d(655) xor d(654) xor d(650) xor d(648) xor d(647) xor d(642) xor d(640) xor d(637) xor d(636) xor d(631) xor d(630) xor d(629) xor d(627) xor d(626) xor d(621) xor d(619) xor d(617) xor d(615) xor d(613) xor d(612) xor d(611) xor d(608) xor d(606) xor d(605) xor d(602) xor d(601) xor d(600) xor d(599) xor d(595) xor d(592) xor d(591) xor d(590) xor d(586) xor d(583) xor d(581) xor d(580) xor d(579) xor d(578) xor d(577) xor d(575) xor d(573) xor d(569) xor d(568) xor d(567) xor d(565) xor d(564) xor d(563) xor d(561) xor d(558) xor d(557) xor d(556) xor d(553) xor d(551) xor d(550) xor d(549) xor d(548) xor d(547) xor d(546) xor d(545) xor d(544) xor d(541) xor d(540) xor d(537) xor d(536) xor d(535) xor d(534) xor d(531) xor d(530) xor d(528) xor d(526) xor d(524) xor d(523) xor d(519) xor d(517) xor d(510) xor d(508) xor d(507) xor d(506) xor d(505) xor d(503) xor d(502) xor d(500) xor d(498) xor d(497) xor d(496) xor d(495) xor d(494) xor d(490) xor d(487) xor d(484) xor d(483) xor d(480) xor d(476) xor d(475) xor d(473) xor d(467) xor d(460) xor d(459) xor d(458) xor d(456) xor d(455) xor d(453) xor d(450) xor d(445) xor d(442) xor d(441) xor d(440) xor d(438) xor d(437) xor d(434) xor d(433) xor d(432) xor d(430) xor d(428) xor d(425) xor d(424) xor d(422) xor d(421) xor d(417) xor d(416) xor d(415) xor d(414) xor d(413) xor d(412) xor d(411) xor d(409) xor d(408) xor d(407) xor d(406) xor d(405) xor d(397) xor d(396) xor d(394) xor d(393) xor d(390) xor d(388) xor d(387) xor d(385) xor d(384) xor d(383) xor d(382) xor d(380) xor d(379) xor d(372) xor d(370) xor d(368) xor d(365) xor d(364) xor d(362) xor d(358) xor d(356) xor d(354) xor d(350) xor d(349) xor d(348) xor d(344) xor d(343) xor d(342) xor d(341) xor d(339) xor d(338) xor d(337) xor d(336) xor d(331) xor d(330) xor d(328) xor d(325) xor d(322) xor d(321) xor d(320) xor d(317) xor d(308) xor d(306) xor d(304) xor d(303) xor d(302) xor d(301) xor d(300) xor d(299) xor d(298) xor d(297) xor d(293) xor d(291) xor d(289) xor d(288) xor d(287) xor d(285) xor d(283) xor d(282) xor d(277) xor d(275) xor d(271) xor d(269) xor d(265) xor d(264) xor d(261) xor d(251) xor d(250) xor d(248) xor d(247) xor d(246) xor d(244) xor d(240) xor d(239) xor d(238) xor d(234) xor d(233) xor d(232) xor d(231) xor d(229) xor d(228) xor d(224) xor d(223) xor d(222) xor d(221) xor d(220) xor d(219) xor d(217) xor d(213) xor d(212) xor d(210) xor d(208) xor d(206) xor d(203) xor d(201) xor d(200) xor d(197) xor d(194) xor d(191) xor d(190) xor d(187) xor d(186) xor d(185) xor d(184) xor d(183) xor d(182) xor d(180) xor d(175) xor d(174) xor d(171) xor d(168) xor d(161) xor d(158) xor d(157) xor d(156) xor d(154) xor d(152) xor d(146) xor d(145) xor d(144) xor d(142) xor d(141) xor d(139) xor d(137) xor d(136) xor d(135) xor d(132) xor d(129) xor d(128) xor d(125) xor d(122) xor d(121) xor d(120) xor d(119) xor d(117) xor d(116) xor d(113) xor d(112) xor d(111) xor d(110) xor d(106) xor d(105) xor d(104) xor d(103) xor d(101) xor d(100) xor d(98) xor d(95) xor d(92) xor d(91) xor d(90) xor d(88) xor d(87) xor d(85) xor d(84) xor d(83) xor d(79) xor d(78) xor d(76) xor d(69) xor d(67) xor d(58) xor d(57) xor d(52) xor d(49) xor d(48) xor d(47) xor d(45) xor d(38) xor d(36) xor d(33) xor d(31) xor d(30) xor d(27) xor d(25) xor d(23) xor d(22) xor d(20) xor d(18) xor d(14) xor d(13) xor d(9) xor d(6) xor d(5) xor d(1) xor c(0) xor c(1) xor c(2) xor c(6) xor c(7) xor c(13) xor c(17) xor c(19) xor c(21) xor c(23) xor c(24) xor c(25) xor c(27) xor c(29) xor c(30) xor c(31);
    newcrc(18) := d(1023) xor d(1022) xor d(1020) xor d(1018) xor d(1017) xor d(1016) xor d(1014) xor d(1012) xor d(1010) xor d(1006) xor d(1000) xor d(999) xor d(995) xor d(994) xor d(993) xor d(992) xor d(991) xor d(990) xor d(989) xor d(987) xor d(986) xor d(981) xor d(980) xor d(978) xor d(977) xor d(975) xor d(974) xor d(973) xor d(971) xor d(969) xor d(968) xor d(967) xor d(966) xor d(965) xor d(964) xor d(963) xor d(962) xor d(961) xor d(960) xor d(959) xor d(957) xor d(956) xor d(952) xor d(950) xor d(948) xor d(947) xor d(946) xor d(945) xor d(943) xor d(942) xor d(941) xor d(940) xor d(937) xor d(936) xor d(935) xor d(934) xor d(928) xor d(927) xor d(924) xor d(923) xor d(921) xor d(920) xor d(919) xor d(917) xor d(916) xor d(915) xor d(914) xor d(911) xor d(909) xor d(907) xor d(905) xor d(904) xor d(902) xor d(900) xor d(899) xor d(898) xor d(895) xor d(894) xor d(889) xor d(888) xor d(886) xor d(883) xor d(879) xor d(875) xor d(872) xor d(871) xor d(870) xor d(867) xor d(865) xor d(864) xor d(859) xor d(858) xor d(853) xor d(851) xor d(850) xor d(848) xor d(843) xor d(839) xor d(835) xor d(834) xor d(833) xor d(832) xor d(825) xor d(824) xor d(822) xor d(820) xor d(818) xor d(817) xor d(816) xor d(815) xor d(812) xor d(808) xor d(807) xor d(806) xor d(803) xor d(801) xor d(800) xor d(796) xor d(795) xor d(794) xor d(787) xor d(785) xor d(782) xor d(780) xor d(777) xor d(775) xor d(772) xor d(769) xor d(765) xor d(764) xor d(763) xor d(752) xor d(751) xor d(748) xor d(747) xor d(746) xor d(742) xor d(741) xor d(739) xor d(738) xor d(735) xor d(731) xor d(730) xor d(728) xor d(727) xor d(725) xor d(719) xor d(718) xor d(716) xor d(712) xor d(711) xor d(709) xor d(708) xor d(704) xor d(701) xor d(698) xor d(695) xor d(694) xor d(693) xor d(692) xor d(691) xor d(687) xor d(686) xor d(681) xor d(680) xor d(678) xor d(677) xor d(676) xor d(673) xor d(671) xor d(666) xor d(665) xor d(664) xor d(662) xor d(660) xor d(657) xor d(656) xor d(655) xor d(651) xor d(649) xor d(648) xor d(643) xor d(641) xor d(638) xor d(637) xor d(632) xor d(631) xor d(630) xor d(628) xor d(627) xor d(622) xor d(620) xor d(618) xor d(616) xor d(614) xor d(613) xor d(612) xor d(609) xor d(607) xor d(606) xor d(603) xor d(602) xor d(601) xor d(600) xor d(596) xor d(593) xor d(592) xor d(591) xor d(587) xor d(584) xor d(582) xor d(581) xor d(580) xor d(579) xor d(578) xor d(576) xor d(574) xor d(570) xor d(569) xor d(568) xor d(566) xor d(565) xor d(564) xor d(562) xor d(559) xor d(558) xor d(557) xor d(554) xor d(552) xor d(551) xor d(550) xor d(549) xor d(548) xor d(547) xor d(546) xor d(545) xor d(542) xor d(541) xor d(538) xor d(537) xor d(536) xor d(535) xor d(532) xor d(531) xor d(529) xor d(527) xor d(525) xor d(524) xor d(520) xor d(518) xor d(511) xor d(509) xor d(508) xor d(507) xor d(506) xor d(504) xor d(503) xor d(501) xor d(499) xor d(498) xor d(497) xor d(496) xor d(495) xor d(491) xor d(488) xor d(485) xor d(484) xor d(481) xor d(477) xor d(476) xor d(474) xor d(468) xor d(461) xor d(460) xor d(459) xor d(457) xor d(456) xor d(454) xor d(451) xor d(446) xor d(443) xor d(442) xor d(441) xor d(439) xor d(438) xor d(435) xor d(434) xor d(433) xor d(431) xor d(429) xor d(426) xor d(425) xor d(423) xor d(422) xor d(418) xor d(417) xor d(416) xor d(415) xor d(414) xor d(413) xor d(412) xor d(410) xor d(409) xor d(408) xor d(407) xor d(406) xor d(398) xor d(397) xor d(395) xor d(394) xor d(391) xor d(389) xor d(388) xor d(386) xor d(385) xor d(384) xor d(383) xor d(381) xor d(380) xor d(373) xor d(371) xor d(369) xor d(366) xor d(365) xor d(363) xor d(359) xor d(357) xor d(355) xor d(351) xor d(350) xor d(349) xor d(345) xor d(344) xor d(343) xor d(342) xor d(340) xor d(339) xor d(338) xor d(337) xor d(332) xor d(331) xor d(329) xor d(326) xor d(323) xor d(322) xor d(321) xor d(318) xor d(309) xor d(307) xor d(305) xor d(304) xor d(303) xor d(302) xor d(301) xor d(300) xor d(299) xor d(298) xor d(294) xor d(292) xor d(290) xor d(289) xor d(288) xor d(286) xor d(284) xor d(283) xor d(278) xor d(276) xor d(272) xor d(270) xor d(266) xor d(265) xor d(262) xor d(252) xor d(251) xor d(249) xor d(248) xor d(247) xor d(245) xor d(241) xor d(240) xor d(239) xor d(235) xor d(234) xor d(233) xor d(232) xor d(230) xor d(229) xor d(225) xor d(224) xor d(223) xor d(222) xor d(221) xor d(220) xor d(218) xor d(214) xor d(213) xor d(211) xor d(209) xor d(207) xor d(204) xor d(202) xor d(201) xor d(198) xor d(195) xor d(192) xor d(191) xor d(188) xor d(187) xor d(186) xor d(185) xor d(184) xor d(183) xor d(181) xor d(176) xor d(175) xor d(172) xor d(169) xor d(162) xor d(159) xor d(158) xor d(157) xor d(155) xor d(153) xor d(147) xor d(146) xor d(145) xor d(143) xor d(142) xor d(140) xor d(138) xor d(137) xor d(136) xor d(133) xor d(130) xor d(129) xor d(126) xor d(123) xor d(122) xor d(121) xor d(120) xor d(118) xor d(117) xor d(114) xor d(113) xor d(112) xor d(111) xor d(107) xor d(106) xor d(105) xor d(104) xor d(102) xor d(101) xor d(99) xor d(96) xor d(93) xor d(92) xor d(91) xor d(89) xor d(88) xor d(86) xor d(85) xor d(84) xor d(80) xor d(79) xor d(77) xor d(70) xor d(68) xor d(59) xor d(58) xor d(53) xor d(50) xor d(49) xor d(48) xor d(46) xor d(39) xor d(37) xor d(34) xor d(32) xor d(31) xor d(28) xor d(26) xor d(24) xor d(23) xor d(21) xor d(19) xor d(15) xor d(14) xor d(10) xor d(7) xor d(6) xor d(2) xor c(0) xor c(1) xor c(2) xor c(3) xor c(7) xor c(8) xor c(14) xor c(18) xor c(20) xor c(22) xor c(24) xor c(25) xor c(26) xor c(28) xor c(30) xor c(31);
    newcrc(19) := d(1023) xor d(1021) xor d(1019) xor d(1018) xor d(1017) xor d(1015) xor d(1013) xor d(1011) xor d(1007) xor d(1001) xor d(1000) xor d(996) xor d(995) xor d(994) xor d(993) xor d(992) xor d(991) xor d(990) xor d(988) xor d(987) xor d(982) xor d(981) xor d(979) xor d(978) xor d(976) xor d(975) xor d(974) xor d(972) xor d(970) xor d(969) xor d(968) xor d(967) xor d(966) xor d(965) xor d(964) xor d(963) xor d(962) xor d(961) xor d(960) xor d(958) xor d(957) xor d(953) xor d(951) xor d(949) xor d(948) xor d(947) xor d(946) xor d(944) xor d(943) xor d(942) xor d(941) xor d(938) xor d(937) xor d(936) xor d(935) xor d(929) xor d(928) xor d(925) xor d(924) xor d(922) xor d(921) xor d(920) xor d(918) xor d(917) xor d(916) xor d(915) xor d(912) xor d(910) xor d(908) xor d(906) xor d(905) xor d(903) xor d(901) xor d(900) xor d(899) xor d(896) xor d(895) xor d(890) xor d(889) xor d(887) xor d(884) xor d(880) xor d(876) xor d(873) xor d(872) xor d(871) xor d(868) xor d(866) xor d(865) xor d(860) xor d(859) xor d(854) xor d(852) xor d(851) xor d(849) xor d(844) xor d(840) xor d(836) xor d(835) xor d(834) xor d(833) xor d(826) xor d(825) xor d(823) xor d(821) xor d(819) xor d(818) xor d(817) xor d(816) xor d(813) xor d(809) xor d(808) xor d(807) xor d(804) xor d(802) xor d(801) xor d(797) xor d(796) xor d(795) xor d(788) xor d(786) xor d(783) xor d(781) xor d(778) xor d(776) xor d(773) xor d(770) xor d(766) xor d(765) xor d(764) xor d(753) xor d(752) xor d(749) xor d(748) xor d(747) xor d(743) xor d(742) xor d(740) xor d(739) xor d(736) xor d(732) xor d(731) xor d(729) xor d(728) xor d(726) xor d(720) xor d(719) xor d(717) xor d(713) xor d(712) xor d(710) xor d(709) xor d(705) xor d(702) xor d(699) xor d(696) xor d(695) xor d(694) xor d(693) xor d(692) xor d(688) xor d(687) xor d(682) xor d(681) xor d(679) xor d(678) xor d(677) xor d(674) xor d(672) xor d(667) xor d(666) xor d(665) xor d(663) xor d(661) xor d(658) xor d(657) xor d(656) xor d(652) xor d(650) xor d(649) xor d(644) xor d(642) xor d(639) xor d(638) xor d(633) xor d(632) xor d(631) xor d(629) xor d(628) xor d(623) xor d(621) xor d(619) xor d(617) xor d(615) xor d(614) xor d(613) xor d(610) xor d(608) xor d(607) xor d(604) xor d(603) xor d(602) xor d(601) xor d(597) xor d(594) xor d(593) xor d(592) xor d(588) xor d(585) xor d(583) xor d(582) xor d(581) xor d(580) xor d(579) xor d(577) xor d(575) xor d(571) xor d(570) xor d(569) xor d(567) xor d(566) xor d(565) xor d(563) xor d(560) xor d(559) xor d(558) xor d(555) xor d(553) xor d(552) xor d(551) xor d(550) xor d(549) xor d(548) xor d(547) xor d(546) xor d(543) xor d(542) xor d(539) xor d(538) xor d(537) xor d(536) xor d(533) xor d(532) xor d(530) xor d(528) xor d(526) xor d(525) xor d(521) xor d(519) xor d(512) xor d(510) xor d(509) xor d(508) xor d(507) xor d(505) xor d(504) xor d(502) xor d(500) xor d(499) xor d(498) xor d(497) xor d(496) xor d(492) xor d(489) xor d(486) xor d(485) xor d(482) xor d(478) xor d(477) xor d(475) xor d(469) xor d(462) xor d(461) xor d(460) xor d(458) xor d(457) xor d(455) xor d(452) xor d(447) xor d(444) xor d(443) xor d(442) xor d(440) xor d(439) xor d(436) xor d(435) xor d(434) xor d(432) xor d(430) xor d(427) xor d(426) xor d(424) xor d(423) xor d(419) xor d(418) xor d(417) xor d(416) xor d(415) xor d(414) xor d(413) xor d(411) xor d(410) xor d(409) xor d(408) xor d(407) xor d(399) xor d(398) xor d(396) xor d(395) xor d(392) xor d(390) xor d(389) xor d(387) xor d(386) xor d(385) xor d(384) xor d(382) xor d(381) xor d(374) xor d(372) xor d(370) xor d(367) xor d(366) xor d(364) xor d(360) xor d(358) xor d(356) xor d(352) xor d(351) xor d(350) xor d(346) xor d(345) xor d(344) xor d(343) xor d(341) xor d(340) xor d(339) xor d(338) xor d(333) xor d(332) xor d(330) xor d(327) xor d(324) xor d(323) xor d(322) xor d(319) xor d(310) xor d(308) xor d(306) xor d(305) xor d(304) xor d(303) xor d(302) xor d(301) xor d(300) xor d(299) xor d(295) xor d(293) xor d(291) xor d(290) xor d(289) xor d(287) xor d(285) xor d(284) xor d(279) xor d(277) xor d(273) xor d(271) xor d(267) xor d(266) xor d(263) xor d(253) xor d(252) xor d(250) xor d(249) xor d(248) xor d(246) xor d(242) xor d(241) xor d(240) xor d(236) xor d(235) xor d(234) xor d(233) xor d(231) xor d(230) xor d(226) xor d(225) xor d(224) xor d(223) xor d(222) xor d(221) xor d(219) xor d(215) xor d(214) xor d(212) xor d(210) xor d(208) xor d(205) xor d(203) xor d(202) xor d(199) xor d(196) xor d(193) xor d(192) xor d(189) xor d(188) xor d(187) xor d(186) xor d(185) xor d(184) xor d(182) xor d(177) xor d(176) xor d(173) xor d(170) xor d(163) xor d(160) xor d(159) xor d(158) xor d(156) xor d(154) xor d(148) xor d(147) xor d(146) xor d(144) xor d(143) xor d(141) xor d(139) xor d(138) xor d(137) xor d(134) xor d(131) xor d(130) xor d(127) xor d(124) xor d(123) xor d(122) xor d(121) xor d(119) xor d(118) xor d(115) xor d(114) xor d(113) xor d(112) xor d(108) xor d(107) xor d(106) xor d(105) xor d(103) xor d(102) xor d(100) xor d(97) xor d(94) xor d(93) xor d(92) xor d(90) xor d(89) xor d(87) xor d(86) xor d(85) xor d(81) xor d(80) xor d(78) xor d(71) xor d(69) xor d(60) xor d(59) xor d(54) xor d(51) xor d(50) xor d(49) xor d(47) xor d(40) xor d(38) xor d(35) xor d(33) xor d(32) xor d(29) xor d(27) xor d(25) xor d(24) xor d(22) xor d(20) xor d(16) xor d(15) xor d(11) xor d(8) xor d(7) xor d(3) xor c(0) xor c(1) xor c(2) xor c(3) xor c(4) xor c(8) xor c(9) xor c(15) xor c(19) xor c(21) xor c(23) xor c(25) xor c(26) xor c(27) xor c(29) xor c(31);
    newcrc(20) := d(1022) xor d(1020) xor d(1019) xor d(1018) xor d(1016) xor d(1014) xor d(1012) xor d(1008) xor d(1002) xor d(1001) xor d(997) xor d(996) xor d(995) xor d(994) xor d(993) xor d(992) xor d(991) xor d(989) xor d(988) xor d(983) xor d(982) xor d(980) xor d(979) xor d(977) xor d(976) xor d(975) xor d(973) xor d(971) xor d(970) xor d(969) xor d(968) xor d(967) xor d(966) xor d(965) xor d(964) xor d(963) xor d(962) xor d(961) xor d(959) xor d(958) xor d(954) xor d(952) xor d(950) xor d(949) xor d(948) xor d(947) xor d(945) xor d(944) xor d(943) xor d(942) xor d(939) xor d(938) xor d(937) xor d(936) xor d(930) xor d(929) xor d(926) xor d(925) xor d(923) xor d(922) xor d(921) xor d(919) xor d(918) xor d(917) xor d(916) xor d(913) xor d(911) xor d(909) xor d(907) xor d(906) xor d(904) xor d(902) xor d(901) xor d(900) xor d(897) xor d(896) xor d(891) xor d(890) xor d(888) xor d(885) xor d(881) xor d(877) xor d(874) xor d(873) xor d(872) xor d(869) xor d(867) xor d(866) xor d(861) xor d(860) xor d(855) xor d(853) xor d(852) xor d(850) xor d(845) xor d(841) xor d(837) xor d(836) xor d(835) xor d(834) xor d(827) xor d(826) xor d(824) xor d(822) xor d(820) xor d(819) xor d(818) xor d(817) xor d(814) xor d(810) xor d(809) xor d(808) xor d(805) xor d(803) xor d(802) xor d(798) xor d(797) xor d(796) xor d(789) xor d(787) xor d(784) xor d(782) xor d(779) xor d(777) xor d(774) xor d(771) xor d(767) xor d(766) xor d(765) xor d(754) xor d(753) xor d(750) xor d(749) xor d(748) xor d(744) xor d(743) xor d(741) xor d(740) xor d(737) xor d(733) xor d(732) xor d(730) xor d(729) xor d(727) xor d(721) xor d(720) xor d(718) xor d(714) xor d(713) xor d(711) xor d(710) xor d(706) xor d(703) xor d(700) xor d(697) xor d(696) xor d(695) xor d(694) xor d(693) xor d(689) xor d(688) xor d(683) xor d(682) xor d(680) xor d(679) xor d(678) xor d(675) xor d(673) xor d(668) xor d(667) xor d(666) xor d(664) xor d(662) xor d(659) xor d(658) xor d(657) xor d(653) xor d(651) xor d(650) xor d(645) xor d(643) xor d(640) xor d(639) xor d(634) xor d(633) xor d(632) xor d(630) xor d(629) xor d(624) xor d(622) xor d(620) xor d(618) xor d(616) xor d(615) xor d(614) xor d(611) xor d(609) xor d(608) xor d(605) xor d(604) xor d(603) xor d(602) xor d(598) xor d(595) xor d(594) xor d(593) xor d(589) xor d(586) xor d(584) xor d(583) xor d(582) xor d(581) xor d(580) xor d(578) xor d(576) xor d(572) xor d(571) xor d(570) xor d(568) xor d(567) xor d(566) xor d(564) xor d(561) xor d(560) xor d(559) xor d(556) xor d(554) xor d(553) xor d(552) xor d(551) xor d(550) xor d(549) xor d(548) xor d(547) xor d(544) xor d(543) xor d(540) xor d(539) xor d(538) xor d(537) xor d(534) xor d(533) xor d(531) xor d(529) xor d(527) xor d(526) xor d(522) xor d(520) xor d(513) xor d(511) xor d(510) xor d(509) xor d(508) xor d(506) xor d(505) xor d(503) xor d(501) xor d(500) xor d(499) xor d(498) xor d(497) xor d(493) xor d(490) xor d(487) xor d(486) xor d(483) xor d(479) xor d(478) xor d(476) xor d(470) xor d(463) xor d(462) xor d(461) xor d(459) xor d(458) xor d(456) xor d(453) xor d(448) xor d(445) xor d(444) xor d(443) xor d(441) xor d(440) xor d(437) xor d(436) xor d(435) xor d(433) xor d(431) xor d(428) xor d(427) xor d(425) xor d(424) xor d(420) xor d(419) xor d(418) xor d(417) xor d(416) xor d(415) xor d(414) xor d(412) xor d(411) xor d(410) xor d(409) xor d(408) xor d(400) xor d(399) xor d(397) xor d(396) xor d(393) xor d(391) xor d(390) xor d(388) xor d(387) xor d(386) xor d(385) xor d(383) xor d(382) xor d(375) xor d(373) xor d(371) xor d(368) xor d(367) xor d(365) xor d(361) xor d(359) xor d(357) xor d(353) xor d(352) xor d(351) xor d(347) xor d(346) xor d(345) xor d(344) xor d(342) xor d(341) xor d(340) xor d(339) xor d(334) xor d(333) xor d(331) xor d(328) xor d(325) xor d(324) xor d(323) xor d(320) xor d(311) xor d(309) xor d(307) xor d(306) xor d(305) xor d(304) xor d(303) xor d(302) xor d(301) xor d(300) xor d(296) xor d(294) xor d(292) xor d(291) xor d(290) xor d(288) xor d(286) xor d(285) xor d(280) xor d(278) xor d(274) xor d(272) xor d(268) xor d(267) xor d(264) xor d(254) xor d(253) xor d(251) xor d(250) xor d(249) xor d(247) xor d(243) xor d(242) xor d(241) xor d(237) xor d(236) xor d(235) xor d(234) xor d(232) xor d(231) xor d(227) xor d(226) xor d(225) xor d(224) xor d(223) xor d(222) xor d(220) xor d(216) xor d(215) xor d(213) xor d(211) xor d(209) xor d(206) xor d(204) xor d(203) xor d(200) xor d(197) xor d(194) xor d(193) xor d(190) xor d(189) xor d(188) xor d(187) xor d(186) xor d(185) xor d(183) xor d(178) xor d(177) xor d(174) xor d(171) xor d(164) xor d(161) xor d(160) xor d(159) xor d(157) xor d(155) xor d(149) xor d(148) xor d(147) xor d(145) xor d(144) xor d(142) xor d(140) xor d(139) xor d(138) xor d(135) xor d(132) xor d(131) xor d(128) xor d(125) xor d(124) xor d(123) xor d(122) xor d(120) xor d(119) xor d(116) xor d(115) xor d(114) xor d(113) xor d(109) xor d(108) xor d(107) xor d(106) xor d(104) xor d(103) xor d(101) xor d(98) xor d(95) xor d(94) xor d(93) xor d(91) xor d(90) xor d(88) xor d(87) xor d(86) xor d(82) xor d(81) xor d(79) xor d(72) xor d(70) xor d(61) xor d(60) xor d(55) xor d(52) xor d(51) xor d(50) xor d(48) xor d(41) xor d(39) xor d(36) xor d(34) xor d(33) xor d(30) xor d(28) xor d(26) xor d(25) xor d(23) xor d(21) xor d(17) xor d(16) xor d(12) xor d(9) xor d(8) xor d(4) xor c(0) xor c(1) xor c(2) xor c(3) xor c(4) xor c(5) xor c(9) xor c(10) xor c(16) xor c(20) xor c(22) xor c(24) xor c(26) xor c(27) xor c(28) xor c(30);
    newcrc(21) := d(1023) xor d(1021) xor d(1020) xor d(1019) xor d(1017) xor d(1015) xor d(1013) xor d(1009) xor d(1003) xor d(1002) xor d(998) xor d(997) xor d(996) xor d(995) xor d(994) xor d(993) xor d(992) xor d(990) xor d(989) xor d(984) xor d(983) xor d(981) xor d(980) xor d(978) xor d(977) xor d(976) xor d(974) xor d(972) xor d(971) xor d(970) xor d(969) xor d(968) xor d(967) xor d(966) xor d(965) xor d(964) xor d(963) xor d(962) xor d(960) xor d(959) xor d(955) xor d(953) xor d(951) xor d(950) xor d(949) xor d(948) xor d(946) xor d(945) xor d(944) xor d(943) xor d(940) xor d(939) xor d(938) xor d(937) xor d(931) xor d(930) xor d(927) xor d(926) xor d(924) xor d(923) xor d(922) xor d(920) xor d(919) xor d(918) xor d(917) xor d(914) xor d(912) xor d(910) xor d(908) xor d(907) xor d(905) xor d(903) xor d(902) xor d(901) xor d(898) xor d(897) xor d(892) xor d(891) xor d(889) xor d(886) xor d(882) xor d(878) xor d(875) xor d(874) xor d(873) xor d(870) xor d(868) xor d(867) xor d(862) xor d(861) xor d(856) xor d(854) xor d(853) xor d(851) xor d(846) xor d(842) xor d(838) xor d(837) xor d(836) xor d(835) xor d(828) xor d(827) xor d(825) xor d(823) xor d(821) xor d(820) xor d(819) xor d(818) xor d(815) xor d(811) xor d(810) xor d(809) xor d(806) xor d(804) xor d(803) xor d(799) xor d(798) xor d(797) xor d(790) xor d(788) xor d(785) xor d(783) xor d(780) xor d(778) xor d(775) xor d(772) xor d(768) xor d(767) xor d(766) xor d(755) xor d(754) xor d(751) xor d(750) xor d(749) xor d(745) xor d(744) xor d(742) xor d(741) xor d(738) xor d(734) xor d(733) xor d(731) xor d(730) xor d(728) xor d(722) xor d(721) xor d(719) xor d(715) xor d(714) xor d(712) xor d(711) xor d(707) xor d(704) xor d(701) xor d(698) xor d(697) xor d(696) xor d(695) xor d(694) xor d(690) xor d(689) xor d(684) xor d(683) xor d(681) xor d(680) xor d(679) xor d(676) xor d(674) xor d(669) xor d(668) xor d(667) xor d(665) xor d(663) xor d(660) xor d(659) xor d(658) xor d(654) xor d(652) xor d(651) xor d(646) xor d(644) xor d(641) xor d(640) xor d(635) xor d(634) xor d(633) xor d(631) xor d(630) xor d(625) xor d(623) xor d(621) xor d(619) xor d(617) xor d(616) xor d(615) xor d(612) xor d(610) xor d(609) xor d(606) xor d(605) xor d(604) xor d(603) xor d(599) xor d(596) xor d(595) xor d(594) xor d(590) xor d(587) xor d(585) xor d(584) xor d(583) xor d(582) xor d(581) xor d(579) xor d(577) xor d(573) xor d(572) xor d(571) xor d(569) xor d(568) xor d(567) xor d(565) xor d(562) xor d(561) xor d(560) xor d(557) xor d(555) xor d(554) xor d(553) xor d(552) xor d(551) xor d(550) xor d(549) xor d(548) xor d(545) xor d(544) xor d(541) xor d(540) xor d(539) xor d(538) xor d(535) xor d(534) xor d(532) xor d(530) xor d(528) xor d(527) xor d(523) xor d(521) xor d(514) xor d(512) xor d(511) xor d(510) xor d(509) xor d(507) xor d(506) xor d(504) xor d(502) xor d(501) xor d(500) xor d(499) xor d(498) xor d(494) xor d(491) xor d(488) xor d(487) xor d(484) xor d(480) xor d(479) xor d(477) xor d(471) xor d(464) xor d(463) xor d(462) xor d(460) xor d(459) xor d(457) xor d(454) xor d(449) xor d(446) xor d(445) xor d(444) xor d(442) xor d(441) xor d(438) xor d(437) xor d(436) xor d(434) xor d(432) xor d(429) xor d(428) xor d(426) xor d(425) xor d(421) xor d(420) xor d(419) xor d(418) xor d(417) xor d(416) xor d(415) xor d(413) xor d(412) xor d(411) xor d(410) xor d(409) xor d(401) xor d(400) xor d(398) xor d(397) xor d(394) xor d(392) xor d(391) xor d(389) xor d(388) xor d(387) xor d(386) xor d(384) xor d(383) xor d(376) xor d(374) xor d(372) xor d(369) xor d(368) xor d(366) xor d(362) xor d(360) xor d(358) xor d(354) xor d(353) xor d(352) xor d(348) xor d(347) xor d(346) xor d(345) xor d(343) xor d(342) xor d(341) xor d(340) xor d(335) xor d(334) xor d(332) xor d(329) xor d(326) xor d(325) xor d(324) xor d(321) xor d(312) xor d(310) xor d(308) xor d(307) xor d(306) xor d(305) xor d(304) xor d(303) xor d(302) xor d(301) xor d(297) xor d(295) xor d(293) xor d(292) xor d(291) xor d(289) xor d(287) xor d(286) xor d(281) xor d(279) xor d(275) xor d(273) xor d(269) xor d(268) xor d(265) xor d(255) xor d(254) xor d(252) xor d(251) xor d(250) xor d(248) xor d(244) xor d(243) xor d(242) xor d(238) xor d(237) xor d(236) xor d(235) xor d(233) xor d(232) xor d(228) xor d(227) xor d(226) xor d(225) xor d(224) xor d(223) xor d(221) xor d(217) xor d(216) xor d(214) xor d(212) xor d(210) xor d(207) xor d(205) xor d(204) xor d(201) xor d(198) xor d(195) xor d(194) xor d(191) xor d(190) xor d(189) xor d(188) xor d(187) xor d(186) xor d(184) xor d(179) xor d(178) xor d(175) xor d(172) xor d(165) xor d(162) xor d(161) xor d(160) xor d(158) xor d(156) xor d(150) xor d(149) xor d(148) xor d(146) xor d(145) xor d(143) xor d(141) xor d(140) xor d(139) xor d(136) xor d(133) xor d(132) xor d(129) xor d(126) xor d(125) xor d(124) xor d(123) xor d(121) xor d(120) xor d(117) xor d(116) xor d(115) xor d(114) xor d(110) xor d(109) xor d(108) xor d(107) xor d(105) xor d(104) xor d(102) xor d(99) xor d(96) xor d(95) xor d(94) xor d(92) xor d(91) xor d(89) xor d(88) xor d(87) xor d(83) xor d(82) xor d(80) xor d(73) xor d(71) xor d(62) xor d(61) xor d(56) xor d(53) xor d(52) xor d(51) xor d(49) xor d(42) xor d(40) xor d(37) xor d(35) xor d(34) xor d(31) xor d(29) xor d(27) xor d(26) xor d(24) xor d(22) xor d(18) xor d(17) xor d(13) xor d(10) xor d(9) xor d(5) xor c(0) xor c(1) xor c(2) xor c(3) xor c(4) xor c(5) xor c(6) xor c(10) xor c(11) xor c(17) xor c(21) xor c(23) xor c(25) xor c(27) xor c(28) xor c(29) xor c(31);
    newcrc(22) := d(1022) xor d(1020) xor d(1019) xor d(1015) xor d(1014) xor d(1012) xor d(1011) xor d(1010) xor d(1009) xor d(1008) xor d(1006) xor d(1005) xor d(1003) xor d(1000) xor d(997) xor d(995) xor d(993) xor d(992) xor d(991) xor d(983) xor d(980) xor d(974) xor d(973) xor d(972) xor d(970) xor d(969) xor d(968) xor d(966) xor d(965) xor d(964) xor d(963) xor d(961) xor d(959) xor d(958) xor d(956) xor d(955) xor d(953) xor d(952) xor d(951) xor d(949) xor d(948) xor d(947) xor d(946) xor d(945) xor d(940) xor d(935) xor d(934) xor d(933) xor d(932) xor d(928) xor d(927) xor d(925) xor d(924) xor d(923) xor d(921) xor d(919) xor d(917) xor d(913) xor d(911) xor d(910) xor d(909) xor d(908) xor d(907) xor d(901) xor d(900) xor d(897) xor d(896) xor d(892) xor d(891) xor d(889) xor d(886) xor d(881) xor d(878) xor d(877) xor d(873) xor d(867) xor d(862) xor d(861) xor d(860) xor d(859) xor d(855) xor d(853) xor d(852) xor d(851) xor d(850) xor d(849) xor d(848) xor d(847) xor d(846) xor d(843) xor d(842) xor d(840) xor d(838) xor d(836) xor d(835) xor d(834) xor d(832) xor d(829) xor d(828) xor d(827) xor d(826) xor d(825) xor d(822) xor d(821) xor d(820) xor d(818) xor d(815) xor d(814) xor d(813) xor d(809) xor d(808) xor d(806) xor d(805) xor d(803) xor d(802) xor d(799) xor d(793) xor d(789) xor d(788) xor d(785) xor d(782) xor d(781) xor d(780) xor d(779) xor d(774) xor d(773) xor d(768) xor d(765) xor d(763) xor d(762) xor d(758) xor d(753) xor d(752) xor d(751) xor d(748) xor d(747) xor d(746) xor d(745) xor d(744) xor d(743) xor d(741) xor d(740) xor d(739) xor d(736) xor d(735) xor d(734) xor d(727) xor d(725) xor d(724) xor d(721) xor d(719) xor d(716) xor d(713) xor d(712) xor d(710) xor d(707) xor d(705) xor d(704) xor d(701) xor d(700) xor d(699) xor d(697) xor d(696) xor d(694) xor d(693) xor d(690) xor d(689) xor d(687) xor d(686) xor d(685) xor d(684) xor d(682) xor d(681) xor d(677) xor d(674) xor d(673) xor d(672) xor d(667) xor d(665) xor d(664) xor d(661) xor d(660) xor d(659) xor d(658) xor d(656) xor d(649) xor d(648) xor d(647) xor d(646) xor d(645) xor d(644) xor d(641) xor d(640) xor d(635) xor d(634) xor d(631) xor d(630) xor d(629) xor d(623) xor d(622) xor d(619) xor d(618) xor d(616) xor d(615) xor d(612) xor d(609) xor d(605) xor d(603) xor d(602) xor d(599) xor d(597) xor d(593) xor d(592) xor d(588) xor d(587) xor d(584) xor d(582) xor d(575) xor d(572) xor d(571) xor d(570) xor d(569) xor d(568) xor d(567) xor d(566) xor d(565) xor d(562) xor d(560) xor d(557) xor d(553) xor d(552) xor d(550) xor d(546) xor d(541) xor d(536) xor d(534) xor d(533) xor d(532) xor d(530) xor d(526) xor d(525) xor d(524) xor d(521) xor d(519) xor d(518) xor d(516) xor d(515) xor d(514) xor d(513) xor d(506) xor d(505) xor d(503) xor d(499) xor d(494) xor d(493) xor d(491) xor d(490) xor d(486) xor d(485) xor d(483) xor d(482) xor d(479) xor d(478) xor d(477) xor d(476) xor d(470) xor d(468) xor d(463) xor d(462) xor d(460) xor d(455) xor d(452) xor d(449) xor d(448) xor d(447) xor d(446) xor d(445) xor d(444) xor d(443) xor d(442) xor d(439) xor d(438) xor d(436) xor d(435) xor d(434) xor d(430) xor d(429) xor d(427) xor d(426) xor d(424) xor d(421) xor d(420) xor d(417) xor d(413) xor d(411) xor d(410) xor d(409) xor d(408) xor d(407) xor d(405) xor d(404) xor d(402) xor d(401) xor d(400) xor d(396) xor d(395) xor d(391) xor d(389) xor d(386) xor d(385) xor d(384) xor d(381) xor d(378) xor d(377) xor d(376) xor d(375) xor d(374) xor d(373) xor d(372) xor d(370) xor d(368) xor d(367) xor d(366) xor d(362) xor d(361) xor d(358) xor d(357) xor d(355) xor d(354) xor d(346) xor d(345) xor d(343) xor d(339) xor d(338) xor d(337) xor d(336) xor d(334) xor d(330) xor d(328) xor d(326) xor d(325) xor d(321) xor d(320) xor d(319) xor d(318) xor d(317) xor d(315) xor d(313) xor d(312) xor d(311) xor d(310) xor d(308) xor d(307) xor d(306) xor d(304) xor d(300) xor d(299) xor d(297) xor d(295) xor d(293) xor d(286) xor d(283) xor d(282) xor d(280) xor d(279) xor d(277) xor d(273) xor d(270) xor d(268) xor d(266) xor d(265) xor d(264) xor d(261) xor d(259) xor d(257) xor d(256) xor d(253) xor d(251) xor d(249) xor d(248) xor d(245) xor d(244) xor d(239) xor d(238) xor d(236) xor d(233) xor d(230) xor d(229) xor d(225) xor d(222) xor d(218) xor d(217) xor d(216) xor d(215) xor d(214) xor d(213) xor d(212) xor d(211) xor d(210) xor d(209) xor d(207) xor d(206) xor d(205) xor d(203) xor d(201) xor d(198) xor d(197) xor d(196) xor d(195) xor d(194) xor d(193) xor d(189) xor d(187) xor d(186) xor d(185) xor d(183) xor d(182) xor d(180) xor d(179) xor d(176) xor d(173) xor d(172) xor d(171) xor d(170) xor d(169) xor d(167) xor d(163) xor d(159) xor d(158) xor d(157) xor d(156) xor d(155) xor d(150) xor d(147) xor d(146) xor d(143) xor d(142) xor d(141) xor d(140) xor d(136) xor d(135) xor d(133) xor d(132) xor d(130) xor d(128) xor d(124) xor d(123) xor d(122) xor d(121) xor d(119) xor d(115) xor d(114) xor d(113) xor d(109) xor d(108) xor d(105) xor d(104) xor d(101) xor d(100) xor d(99) xor d(98) xor d(94) xor d(93) xor d(92) xor d(90) xor d(89) xor d(88) xor d(87) xor d(85) xor d(82) xor d(79) xor d(74) xor d(73) xor d(68) xor d(67) xor d(66) xor d(65) xor d(62) xor d(61) xor d(60) xor d(58) xor d(57) xor d(55) xor d(52) xor d(48) xor d(47) xor d(45) xor d(44) xor d(43) xor d(41) xor d(38) xor d(37) xor d(36) xor d(35) xor d(34) xor d(31) xor d(29) xor d(27) xor d(26) xor d(24) xor d(23) xor d(19) xor d(18) xor d(16) xor d(14) xor d(12) xor d(11) xor d(9) xor d(0) xor c(0) xor c(1) xor c(3) xor c(5) xor c(8) xor c(11) xor c(13) xor c(14) xor c(16) xor c(17) xor c(18) xor c(19) xor c(20) xor c(22) xor c(23) xor c(27) xor c(28) xor c(30);
    newcrc(23) := d(1023) xor d(1020) xor d(1019) xor d(1018) xor d(1013) xor d(1010) xor d(1008) xor d(1007) xor d(1005) xor d(1001) xor d(1000) xor d(999) xor d(993) xor d(990) xor d(985) xor d(983) xor d(982) xor d(980) xor d(979) xor d(978) xor d(977) xor d(973) xor d(970) xor d(969) xor d(966) xor d(965) xor d(964) xor d(962) xor d(958) xor d(957) xor d(956) xor d(955) xor d(952) xor d(949) xor d(947) xor d(946) xor d(944) xor d(939) xor d(938) xor d(936) xor d(931) xor d(929) xor d(928) xor d(926) xor d(925) xor d(924) xor d(922) xor d(917) xor d(915) xor d(914) xor d(912) xor d(911) xor d(909) xor d(908) xor d(907) xor d(906) xor d(904) xor d(903) xor d(900) xor d(899) xor d(896) xor d(892) xor d(891) xor d(889) xor d(886) xor d(883) xor d(882) xor d(881) xor d(877) xor d(876) xor d(875) xor d(873) xor d(871) xor d(869) xor d(867) xor d(862) xor d(859) xor d(857) xor d(856) xor d(852) xor d(847) xor d(846) xor d(844) xor d(843) xor d(842) xor d(841) xor d(840) xor d(836) xor d(834) xor d(833) xor d(832) xor d(830) xor d(829) xor d(828) xor d(826) xor d(825) xor d(824) xor d(823) xor d(822) xor d(821) xor d(818) xor d(813) xor d(812) xor d(811) xor d(808) xor d(802) xor d(798) xor d(794) xor d(793) xor d(791) xor d(790) xor d(789) xor d(788) xor d(785) xor d(784) xor d(783) xor d(781) xor d(776) xor d(775) xor d(767) xor d(766) xor d(765) xor d(764) xor d(762) xor d(759) xor d(758) xor d(756) xor d(755) xor d(754) xor d(752) xor d(750) xor d(749) xor d(746) xor d(745) xor d(737) xor d(735) xor d(732) xor d(731) xor d(729) xor d(728) xor d(727) xor d(726) xor d(724) xor d(723) xor d(721) xor d(719) xor d(717) xor d(715) xor d(714) xor d(713) xor d(711) xor d(710) xor d(707) xor d(706) xor d(705) xor d(704) xor d(697) xor d(693) xor d(690) xor d(689) xor d(688) xor d(685) xor d(683) xor d(682) xor d(680) xor d(678) xor d(672) xor d(670) xor d(669) xor d(667) xor d(662) xor d(661) xor d(660) xor d(659) xor d(658) xor d(657) xor d(656) xor d(655) xor d(653) xor d(652) xor d(650) xor d(647) xor d(645) xor d(644) xor d(641) xor d(640) xor d(635) xor d(631) xor d(629) xor d(626) xor d(616) xor d(615) xor d(612) xor d(611) xor d(609) xor d(607) xor d(602) xor d(599) xor d(598) xor d(596) xor d(595) xor d(594) xor d(592) xor d(591) xor d(589) xor d(588) xor d(587) xor d(586) xor d(580) xor d(578) xor d(576) xor d(575) xor d(574) xor d(572) xor d(570) xor d(569) xor d(568) xor d(566) xor d(565) xor d(560) xor d(557) xor d(556) xor d(555) xor d(553) xor d(549) xor d(547) xor d(545) xor d(540) xor d(539) xor d(537) xor d(533) xor d(532) xor d(530) xor d(529) xor d(528) xor d(527) xor d(521) xor d(520) xor d(518) xor d(517) xor d(515) xor d(512) xor d(511) xor d(510) xor d(508) xor d(504) xor d(502) xor d(501) xor d(493) xor d(490) xor d(489) xor d(488) xor d(487) xor d(484) xor d(482) xor d(481) xor d(478) xor d(476) xor d(472) xor d(471) xor d(470) xor d(469) xor d(468) xor d(465) xor d(463) xor d(462) xor d(458) xor d(456) xor d(453) xor d(452) xor d(447) xor d(446) xor d(445) xor d(443) xor d(440) xor d(439) xor d(435) xor d(434) xor d(433) xor d(431) xor d(430) xor d(428) xor d(427) xor d(425) xor d(424) xor d(421) xor d(419) xor d(416) xor d(411) xor d(410) xor d(407) xor d(406) xor d(404) xor d(403) xor d(402) xor d(401) xor d(400) xor d(399) xor d(398) xor d(397) xor d(393) xor d(391) xor d(388) xor d(385) xor d(382) xor d(381) xor d(379) xor d(377) xor d(375) xor d(373) xor d(372) xor d(371) xor d(367) xor d(366) xor d(357) xor d(356) xor d(355) xor d(353) xor d(349) xor d(348) xor d(346) xor d(345) xor d(342) xor d(341) xor d(340) xor d(334) xor d(333) xor d(331) xor d(329) xor d(328) xor d(326) xor d(317) xor d(316) xor d(315) xor d(314) xor d(313) xor d(311) xor d(310) xor d(308) xor d(307) xor d(303) xor d(302) xor d(301) xor d(299) xor d(297) xor d(295) xor d(292) xor d(290) xor d(288) xor d(286) xor d(284) xor d(281) xor d(280) xor d(279) xor d(278) xor d(277) xor d(276) xor d(273) xor d(271) xor d(268) xor d(267) xor d(266) xor d(264) xor d(262) xor d(261) xor d(260) xor d(259) xor d(258) xor d(255) xor d(254) xor d(250) xor d(249) xor d(248) xor d(246) xor d(245) xor d(243) xor d(240) xor d(239) xor d(231) xor d(228) xor d(227) xor d(224) xor d(223) xor d(219) xor d(218) xor d(217) xor d(215) xor d(213) xor d(211) xor d(209) xor d(206) xor d(204) xor d(203) xor d(201) xor d(196) xor d(195) xor d(193) xor d(192) xor d(191) xor d(187) xor d(184) xor d(182) xor d(181) xor d(180) xor d(177) xor d(174) xor d(173) xor d(169) xor d(168) xor d(167) xor d(166) xor d(164) xor d(162) xor d(161) xor d(160) xor d(159) xor d(157) xor d(155) xor d(149) xor d(148) xor d(147) xor d(142) xor d(141) xor d(135) xor d(133) xor d(132) xor d(131) xor d(129) xor d(128) xor d(127) xor d(126) xor d(124) xor d(122) xor d(120) xor d(119) xor d(118) xor d(117) xor d(115) xor d(113) xor d(111) xor d(109) xor d(105) xor d(104) xor d(103) xor d(102) xor d(100) xor d(98) xor d(97) xor d(96) xor d(93) xor d(91) xor d(90) xor d(89) xor d(88) xor d(87) xor d(86) xor d(85) xor d(84) xor d(82) xor d(81) xor d(80) xor d(79) xor d(75) xor d(74) xor d(73) xor d(72) xor d(69) xor d(65) xor d(62) xor d(60) xor d(59) xor d(56) xor d(55) xor d(54) xor d(50) xor d(49) xor d(47) xor d(46) xor d(42) xor d(39) xor d(38) xor d(36) xor d(35) xor d(34) xor d(31) xor d(29) xor d(27) xor d(26) xor d(20) xor d(19) xor d(17) xor d(16) xor d(15) xor d(13) xor d(9) xor d(6) xor d(1) xor d(0) xor c(1) xor c(7) xor c(8) xor c(9) xor c(13) xor c(15) xor c(16) xor c(18) xor c(21) xor c(26) xor c(27) xor c(28) xor c(31);
    newcrc(24) := d(1021) xor d(1020) xor d(1019) xor d(1014) xor d(1011) xor d(1009) xor d(1008) xor d(1006) xor d(1002) xor d(1001) xor d(1000) xor d(994) xor d(991) xor d(986) xor d(984) xor d(983) xor d(981) xor d(980) xor d(979) xor d(978) xor d(974) xor d(971) xor d(970) xor d(967) xor d(966) xor d(965) xor d(963) xor d(959) xor d(958) xor d(957) xor d(956) xor d(953) xor d(950) xor d(948) xor d(947) xor d(945) xor d(940) xor d(939) xor d(937) xor d(932) xor d(930) xor d(929) xor d(927) xor d(926) xor d(925) xor d(923) xor d(918) xor d(916) xor d(915) xor d(913) xor d(912) xor d(910) xor d(909) xor d(908) xor d(907) xor d(905) xor d(904) xor d(901) xor d(900) xor d(897) xor d(893) xor d(892) xor d(890) xor d(887) xor d(884) xor d(883) xor d(882) xor d(878) xor d(877) xor d(876) xor d(874) xor d(872) xor d(870) xor d(868) xor d(863) xor d(860) xor d(858) xor d(857) xor d(853) xor d(848) xor d(847) xor d(845) xor d(844) xor d(843) xor d(842) xor d(841) xor d(837) xor d(835) xor d(834) xor d(833) xor d(831) xor d(830) xor d(829) xor d(827) xor d(826) xor d(825) xor d(824) xor d(823) xor d(822) xor d(819) xor d(814) xor d(813) xor d(812) xor d(809) xor d(803) xor d(799) xor d(795) xor d(794) xor d(792) xor d(791) xor d(790) xor d(789) xor d(786) xor d(785) xor d(784) xor d(782) xor d(777) xor d(776) xor d(768) xor d(767) xor d(766) xor d(765) xor d(763) xor d(760) xor d(759) xor d(757) xor d(756) xor d(755) xor d(753) xor d(751) xor d(750) xor d(747) xor d(746) xor d(738) xor d(736) xor d(733) xor d(732) xor d(730) xor d(729) xor d(728) xor d(727) xor d(725) xor d(724) xor d(722) xor d(720) xor d(718) xor d(716) xor d(715) xor d(714) xor d(712) xor d(711) xor d(708) xor d(707) xor d(706) xor d(705) xor d(698) xor d(694) xor d(691) xor d(690) xor d(689) xor d(686) xor d(684) xor d(683) xor d(681) xor d(679) xor d(673) xor d(671) xor d(670) xor d(668) xor d(663) xor d(662) xor d(661) xor d(660) xor d(659) xor d(658) xor d(657) xor d(656) xor d(654) xor d(653) xor d(651) xor d(648) xor d(646) xor d(645) xor d(642) xor d(641) xor d(636) xor d(632) xor d(630) xor d(627) xor d(617) xor d(616) xor d(613) xor d(612) xor d(610) xor d(608) xor d(603) xor d(600) xor d(599) xor d(597) xor d(596) xor d(595) xor d(593) xor d(592) xor d(590) xor d(589) xor d(588) xor d(587) xor d(581) xor d(579) xor d(577) xor d(576) xor d(575) xor d(573) xor d(571) xor d(570) xor d(569) xor d(567) xor d(566) xor d(561) xor d(558) xor d(557) xor d(556) xor d(554) xor d(550) xor d(548) xor d(546) xor d(541) xor d(540) xor d(538) xor d(534) xor d(533) xor d(531) xor d(530) xor d(529) xor d(528) xor d(522) xor d(521) xor d(519) xor d(518) xor d(516) xor d(513) xor d(512) xor d(511) xor d(509) xor d(505) xor d(503) xor d(502) xor d(494) xor d(491) xor d(490) xor d(489) xor d(488) xor d(485) xor d(483) xor d(482) xor d(479) xor d(477) xor d(473) xor d(472) xor d(471) xor d(470) xor d(469) xor d(466) xor d(464) xor d(463) xor d(459) xor d(457) xor d(454) xor d(453) xor d(448) xor d(447) xor d(446) xor d(444) xor d(441) xor d(440) xor d(436) xor d(435) xor d(434) xor d(432) xor d(431) xor d(429) xor d(428) xor d(426) xor d(425) xor d(422) xor d(420) xor d(417) xor d(412) xor d(411) xor d(408) xor d(407) xor d(405) xor d(404) xor d(403) xor d(402) xor d(401) xor d(400) xor d(399) xor d(398) xor d(394) xor d(392) xor d(389) xor d(386) xor d(383) xor d(382) xor d(380) xor d(378) xor d(376) xor d(374) xor d(373) xor d(372) xor d(368) xor d(367) xor d(358) xor d(357) xor d(356) xor d(354) xor d(350) xor d(349) xor d(347) xor d(346) xor d(343) xor d(342) xor d(341) xor d(335) xor d(334) xor d(332) xor d(330) xor d(329) xor d(327) xor d(318) xor d(317) xor d(316) xor d(315) xor d(314) xor d(312) xor d(311) xor d(309) xor d(308) xor d(304) xor d(303) xor d(302) xor d(300) xor d(298) xor d(296) xor d(293) xor d(291) xor d(289) xor d(287) xor d(285) xor d(282) xor d(281) xor d(280) xor d(279) xor d(278) xor d(277) xor d(274) xor d(272) xor d(269) xor d(268) xor d(267) xor d(265) xor d(263) xor d(262) xor d(261) xor d(260) xor d(259) xor d(256) xor d(255) xor d(251) xor d(250) xor d(249) xor d(247) xor d(246) xor d(244) xor d(241) xor d(240) xor d(232) xor d(229) xor d(228) xor d(225) xor d(224) xor d(220) xor d(219) xor d(218) xor d(216) xor d(214) xor d(212) xor d(210) xor d(207) xor d(205) xor d(204) xor d(202) xor d(197) xor d(196) xor d(194) xor d(193) xor d(192) xor d(188) xor d(185) xor d(183) xor d(182) xor d(181) xor d(178) xor d(175) xor d(174) xor d(170) xor d(169) xor d(168) xor d(167) xor d(165) xor d(163) xor d(162) xor d(161) xor d(160) xor d(158) xor d(156) xor d(150) xor d(149) xor d(148) xor d(143) xor d(142) xor d(136) xor d(134) xor d(133) xor d(132) xor d(130) xor d(129) xor d(128) xor d(127) xor d(125) xor d(123) xor d(121) xor d(120) xor d(119) xor d(118) xor d(116) xor d(114) xor d(112) xor d(110) xor d(106) xor d(105) xor d(104) xor d(103) xor d(101) xor d(99) xor d(98) xor d(97) xor d(94) xor d(92) xor d(91) xor d(90) xor d(89) xor d(88) xor d(87) xor d(86) xor d(85) xor d(83) xor d(82) xor d(81) xor d(80) xor d(76) xor d(75) xor d(74) xor d(73) xor d(70) xor d(66) xor d(63) xor d(61) xor d(60) xor d(57) xor d(56) xor d(55) xor d(51) xor d(50) xor d(48) xor d(47) xor d(43) xor d(40) xor d(39) xor d(37) xor d(36) xor d(35) xor d(32) xor d(30) xor d(28) xor d(27) xor d(21) xor d(20) xor d(18) xor d(17) xor d(16) xor d(14) xor d(10) xor d(7) xor d(2) xor d(1) xor c(2) xor c(8) xor c(9) xor c(10) xor c(14) xor c(16) xor c(17) xor c(19) xor c(22) xor c(27) xor c(28) xor c(29);
    newcrc(25) := d(1022) xor d(1021) xor d(1020) xor d(1015) xor d(1012) xor d(1010) xor d(1009) xor d(1007) xor d(1003) xor d(1002) xor d(1001) xor d(995) xor d(992) xor d(987) xor d(985) xor d(984) xor d(982) xor d(981) xor d(980) xor d(979) xor d(975) xor d(972) xor d(971) xor d(968) xor d(967) xor d(966) xor d(964) xor d(960) xor d(959) xor d(958) xor d(957) xor d(954) xor d(951) xor d(949) xor d(948) xor d(946) xor d(941) xor d(940) xor d(938) xor d(933) xor d(931) xor d(930) xor d(928) xor d(927) xor d(926) xor d(924) xor d(919) xor d(917) xor d(916) xor d(914) xor d(913) xor d(911) xor d(910) xor d(909) xor d(908) xor d(906) xor d(905) xor d(902) xor d(901) xor d(898) xor d(894) xor d(893) xor d(891) xor d(888) xor d(885) xor d(884) xor d(883) xor d(879) xor d(878) xor d(877) xor d(875) xor d(873) xor d(871) xor d(869) xor d(864) xor d(861) xor d(859) xor d(858) xor d(854) xor d(849) xor d(848) xor d(846) xor d(845) xor d(844) xor d(843) xor d(842) xor d(838) xor d(836) xor d(835) xor d(834) xor d(832) xor d(831) xor d(830) xor d(828) xor d(827) xor d(826) xor d(825) xor d(824) xor d(823) xor d(820) xor d(815) xor d(814) xor d(813) xor d(810) xor d(804) xor d(800) xor d(796) xor d(795) xor d(793) xor d(792) xor d(791) xor d(790) xor d(787) xor d(786) xor d(785) xor d(783) xor d(778) xor d(777) xor d(769) xor d(768) xor d(767) xor d(766) xor d(764) xor d(761) xor d(760) xor d(758) xor d(757) xor d(756) xor d(754) xor d(752) xor d(751) xor d(748) xor d(747) xor d(739) xor d(737) xor d(734) xor d(733) xor d(731) xor d(730) xor d(729) xor d(728) xor d(726) xor d(725) xor d(723) xor d(721) xor d(719) xor d(717) xor d(716) xor d(715) xor d(713) xor d(712) xor d(709) xor d(708) xor d(707) xor d(706) xor d(699) xor d(695) xor d(692) xor d(691) xor d(690) xor d(687) xor d(685) xor d(684) xor d(682) xor d(680) xor d(674) xor d(672) xor d(671) xor d(669) xor d(664) xor d(663) xor d(662) xor d(661) xor d(660) xor d(659) xor d(658) xor d(657) xor d(655) xor d(654) xor d(652) xor d(649) xor d(647) xor d(646) xor d(643) xor d(642) xor d(637) xor d(633) xor d(631) xor d(628) xor d(618) xor d(617) xor d(614) xor d(613) xor d(611) xor d(609) xor d(604) xor d(601) xor d(600) xor d(598) xor d(597) xor d(596) xor d(594) xor d(593) xor d(591) xor d(590) xor d(589) xor d(588) xor d(582) xor d(580) xor d(578) xor d(577) xor d(576) xor d(574) xor d(572) xor d(571) xor d(570) xor d(568) xor d(567) xor d(562) xor d(559) xor d(558) xor d(557) xor d(555) xor d(551) xor d(549) xor d(547) xor d(542) xor d(541) xor d(539) xor d(535) xor d(534) xor d(532) xor d(531) xor d(530) xor d(529) xor d(523) xor d(522) xor d(520) xor d(519) xor d(517) xor d(514) xor d(513) xor d(512) xor d(510) xor d(506) xor d(504) xor d(503) xor d(495) xor d(492) xor d(491) xor d(490) xor d(489) xor d(486) xor d(484) xor d(483) xor d(480) xor d(478) xor d(474) xor d(473) xor d(472) xor d(471) xor d(470) xor d(467) xor d(465) xor d(464) xor d(460) xor d(458) xor d(455) xor d(454) xor d(449) xor d(448) xor d(447) xor d(445) xor d(442) xor d(441) xor d(437) xor d(436) xor d(435) xor d(433) xor d(432) xor d(430) xor d(429) xor d(427) xor d(426) xor d(423) xor d(421) xor d(418) xor d(413) xor d(412) xor d(409) xor d(408) xor d(406) xor d(405) xor d(404) xor d(403) xor d(402) xor d(401) xor d(400) xor d(399) xor d(395) xor d(393) xor d(390) xor d(387) xor d(384) xor d(383) xor d(381) xor d(379) xor d(377) xor d(375) xor d(374) xor d(373) xor d(369) xor d(368) xor d(359) xor d(358) xor d(357) xor d(355) xor d(351) xor d(350) xor d(348) xor d(347) xor d(344) xor d(343) xor d(342) xor d(336) xor d(335) xor d(333) xor d(331) xor d(330) xor d(328) xor d(319) xor d(318) xor d(317) xor d(316) xor d(315) xor d(313) xor d(312) xor d(310) xor d(309) xor d(305) xor d(304) xor d(303) xor d(301) xor d(299) xor d(297) xor d(294) xor d(292) xor d(290) xor d(288) xor d(286) xor d(283) xor d(282) xor d(281) xor d(280) xor d(279) xor d(278) xor d(275) xor d(273) xor d(270) xor d(269) xor d(268) xor d(266) xor d(264) xor d(263) xor d(262) xor d(261) xor d(260) xor d(257) xor d(256) xor d(252) xor d(251) xor d(250) xor d(248) xor d(247) xor d(245) xor d(242) xor d(241) xor d(233) xor d(230) xor d(229) xor d(226) xor d(225) xor d(221) xor d(220) xor d(219) xor d(217) xor d(215) xor d(213) xor d(211) xor d(208) xor d(206) xor d(205) xor d(203) xor d(198) xor d(197) xor d(195) xor d(194) xor d(193) xor d(189) xor d(186) xor d(184) xor d(183) xor d(182) xor d(179) xor d(176) xor d(175) xor d(171) xor d(170) xor d(169) xor d(168) xor d(166) xor d(164) xor d(163) xor d(162) xor d(161) xor d(159) xor d(157) xor d(151) xor d(150) xor d(149) xor d(144) xor d(143) xor d(137) xor d(135) xor d(134) xor d(133) xor d(131) xor d(130) xor d(129) xor d(128) xor d(126) xor d(124) xor d(122) xor d(121) xor d(120) xor d(119) xor d(117) xor d(115) xor d(113) xor d(111) xor d(107) xor d(106) xor d(105) xor d(104) xor d(102) xor d(100) xor d(99) xor d(98) xor d(95) xor d(93) xor d(92) xor d(91) xor d(90) xor d(89) xor d(88) xor d(87) xor d(86) xor d(84) xor d(83) xor d(82) xor d(81) xor d(77) xor d(76) xor d(75) xor d(74) xor d(71) xor d(67) xor d(64) xor d(62) xor d(61) xor d(58) xor d(57) xor d(56) xor d(52) xor d(51) xor d(49) xor d(48) xor d(44) xor d(41) xor d(40) xor d(38) xor d(37) xor d(36) xor d(33) xor d(31) xor d(29) xor d(28) xor d(22) xor d(21) xor d(19) xor d(18) xor d(17) xor d(15) xor d(11) xor d(8) xor d(3) xor d(2) xor c(0) xor c(3) xor c(9) xor c(10) xor c(11) xor c(15) xor c(17) xor c(18) xor c(20) xor c(23) xor c(28) xor c(29) xor c(30);
    newcrc(26) := d(1023) xor d(1022) xor d(1019) xor d(1018) xor d(1015) xor d(1013) xor d(1012) xor d(1010) xor d(1009) xor d(1006) xor d(1005) xor d(1003) xor d(1002) xor d(1000) xor d(999) xor d(998) xor d(994) xor d(993) xor d(992) xor d(990) xor d(988) xor d(986) xor d(984) xor d(979) xor d(978) xor d(977) xor d(976) xor d(975) xor d(974) xor d(973) xor d(972) xor d(971) xor d(969) xor d(968) xor d(965) xor d(961) xor d(954) xor d(953) xor d(952) xor d(949) xor d(948) xor d(947) xor d(944) xor d(942) xor d(938) xor d(935) xor d(933) xor d(932) xor d(929) xor d(928) xor d(927) xor d(925) xor d(914) xor d(912) xor d(911) xor d(909) xor d(904) xor d(901) xor d(900) xor d(898) xor d(897) xor d(896) xor d(895) xor d(894) xor d(893) xor d(892) xor d(891) xor d(890) xor d(887) xor d(885) xor d(884) xor d(883) xor d(881) xor d(880) xor d(877) xor d(875) xor d(873) xor d(872) xor d(871) xor d(870) xor d(869) xor d(868) xor d(867) xor d(865) xor d(863) xor d(862) xor d(861) xor d(857) xor d(855) xor d(854) xor d(853) xor d(851) xor d(848) xor d(847) xor d(845) xor d(844) xor d(843) xor d(842) xor d(840) xor d(836) xor d(834) xor d(833) xor d(831) xor d(829) xor d(828) xor d(826) xor d(821) xor d(819) xor d(818) xor d(813) xor d(812) xor d(810) xor d(809) xor d(808) xor d(807) xor d(806) xor d(805) xor d(804) xor d(803) xor d(802) xor d(801) xor d(800) xor d(798) xor d(797) xor d(796) xor d(794) xor d(792) xor d(787) xor d(785) xor d(782) xor d(780) xor d(779) xor d(778) xor d(776) xor d(774) xor d(770) xor d(768) xor d(763) xor d(761) xor d(759) xor d(757) xor d(756) xor d(752) xor d(750) xor d(749) xor d(747) xor d(744) xor d(742) xor d(741) xor d(738) xor d(736) xor d(735) xor d(734) xor d(730) xor d(726) xor d(725) xor d(723) xor d(721) xor d(719) xor d(718) xor d(717) xor d(716) xor d(715) xor d(714) xor d(713) xor d(709) xor d(704) xor d(702) xor d(701) xor d(698) xor d(696) xor d(695) xor d(694) xor d(692) xor d(689) xor d(688) xor d(687) xor d(685) xor d(683) xor d(681) xor d(680) xor d(674) xor d(669) xor d(668) xor d(667) xor d(666) xor d(664) xor d(663) xor d(662) xor d(661) xor d(660) xor d(659) xor d(652) xor d(650) xor d(649) xor d(647) xor d(646) xor d(643) xor d(642) xor d(640) xor d(638) xor d(636) xor d(634) xor d(630) xor d(626) xor d(624) xor d(623) xor d(620) xor d(618) xor d(617) xor d(614) xor d(613) xor d(611) xor d(609) xor d(607) xor d(606) xor d(605) xor d(604) xor d(603) xor d(601) xor d(600) xor d(598) xor d(597) xor d(596) xor d(594) xor d(593) xor d(590) xor d(589) xor d(587) xor d(586) xor d(585) xor d(581) xor d(580) xor d(579) xor d(577) xor d(574) xor d(572) xor d(569) xor d(568) xor d(567) xor d(565) xor d(561) xor d(559) xor d(557) xor d(555) xor d(554) xor d(552) xor d(551) xor d(550) xor d(549) xor d(548) xor d(545) xor d(543) xor d(539) xor d(536) xor d(534) xor d(533) xor d(529) xor d(528) xor d(526) xor d(525) xor d(524) xor d(523) xor d(522) xor d(520) xor d(519) xor d(516) xor d(515) xor d(513) xor d(512) xor d(510) xor d(508) xor d(506) xor d(505) xor d(504) xor d(502) xor d(501) xor d(500) xor d(496) xor d(495) xor d(494) xor d(489) xor d(488) xor d(487) xor d(486) xor d(485) xor d(484) xor d(483) xor d(482) xor d(480) xor d(477) xor d(476) xor d(475) xor d(474) xor d(473) xor d(471) xor d(470) xor d(466) xor d(464) xor d(462) xor d(459) xor d(458) xor d(456) xor d(455) xor d(452) xor d(446) xor d(444) xor d(443) xor d(442) xor d(438) xor d(431) xor d(430) xor d(428) xor d(427) xor d(418) xor d(416) xor d(413) xor d(412) xor d(410) xor d(408) xor d(406) xor d(403) xor d(402) xor d(401) xor d(399) xor d(398) xor d(394) xor d(393) xor d(392) xor d(390) xor d(387) xor d(386) xor d(385) xor d(384) xor d(382) xor d(381) xor d(380) xor d(375) xor d(372) xor d(370) xor d(368) xor d(366) xor d(363) xor d(362) xor d(360) xor d(357) xor d(356) xor d(353) xor d(352) xor d(351) xor d(347) xor d(343) xor d(342) xor d(341) xor d(339) xor d(338) xor d(336) xor d(335) xor d(333) xor d(332) xor d(331) xor d(329) xor d(328) xor d(327) xor d(322) xor d(321) xor d(316) xor d(315) xor d(314) xor d(313) xor d(312) xor d(311) xor d(309) xor d(306) xor d(304) xor d(303) xor d(299) xor d(297) xor d(296) xor d(294) xor d(293) xor d(292) xor d(291) xor d(290) xor d(289) xor d(288) xor d(286) xor d(284) xor d(282) xor d(281) xor d(280) xor d(277) xor d(273) xor d(271) xor d(270) xor d(268) xor d(267) xor d(263) xor d(262) xor d(259) xor d(258) xor d(255) xor d(253) xor d(251) xor d(249) xor d(246) xor d(242) xor d(237) xor d(231) xor d(228) xor d(224) xor d(222) xor d(221) xor d(220) xor d(218) xor d(210) xor d(208) xor d(206) xor d(204) xor d(203) xor d(202) xor d(201) xor d(197) xor d(196) xor d(195) xor d(193) xor d(192) xor d(191) xor d(188) xor d(187) xor d(186) xor d(185) xor d(184) xor d(182) xor d(180) xor d(177) xor d(176) xor d(166) xor d(165) xor d(164) xor d(163) xor d(161) xor d(160) xor d(156) xor d(155) xor d(152) xor d(150) xor d(149) xor d(145) xor d(143) xor d(138) xor d(137) xor d(131) xor d(130) xor d(129) xor d(128) xor d(126) xor d(122) xor d(121) xor d(120) xor d(119) xor d(117) xor d(113) xor d(112) xor d(111) xor d(110) xor d(108) xor d(107) xor d(105) xor d(104) xor d(100) xor d(98) xor d(97) xor d(95) xor d(93) xor d(92) xor d(91) xor d(90) xor d(89) xor d(88) xor d(81) xor d(79) xor d(78) xor d(77) xor d(76) xor d(75) xor d(73) xor d(67) xor d(66) xor d(62) xor d(61) xor d(60) xor d(59) xor d(57) xor d(55) xor d(54) xor d(52) xor d(49) xor d(48) xor d(47) xor d(44) xor d(42) xor d(41) xor d(39) xor d(38) xor d(31) xor d(28) xor d(26) xor d(25) xor d(24) xor d(23) xor d(22) xor d(20) xor d(19) xor d(18) xor d(10) xor d(6) xor d(4) xor d(3) xor d(0) xor c(0) xor c(1) xor c(2) xor c(6) xor c(7) xor c(8) xor c(10) xor c(11) xor c(13) xor c(14) xor c(17) xor c(18) xor c(20) xor c(21) xor c(23) xor c(26) xor c(27) xor c(30) xor c(31);
    newcrc(27) := d(1023) xor d(1020) xor d(1019) xor d(1016) xor d(1014) xor d(1013) xor d(1011) xor d(1010) xor d(1007) xor d(1006) xor d(1004) xor d(1003) xor d(1001) xor d(1000) xor d(999) xor d(995) xor d(994) xor d(993) xor d(991) xor d(989) xor d(987) xor d(985) xor d(980) xor d(979) xor d(978) xor d(977) xor d(976) xor d(975) xor d(974) xor d(973) xor d(972) xor d(970) xor d(969) xor d(966) xor d(962) xor d(955) xor d(954) xor d(953) xor d(950) xor d(949) xor d(948) xor d(945) xor d(943) xor d(939) xor d(936) xor d(934) xor d(933) xor d(930) xor d(929) xor d(928) xor d(926) xor d(915) xor d(913) xor d(912) xor d(910) xor d(905) xor d(902) xor d(901) xor d(899) xor d(898) xor d(897) xor d(896) xor d(895) xor d(894) xor d(893) xor d(892) xor d(891) xor d(888) xor d(886) xor d(885) xor d(884) xor d(882) xor d(881) xor d(878) xor d(876) xor d(874) xor d(873) xor d(872) xor d(871) xor d(870) xor d(869) xor d(868) xor d(866) xor d(864) xor d(863) xor d(862) xor d(858) xor d(856) xor d(855) xor d(854) xor d(852) xor d(849) xor d(848) xor d(846) xor d(845) xor d(844) xor d(843) xor d(841) xor d(837) xor d(835) xor d(834) xor d(832) xor d(830) xor d(829) xor d(827) xor d(822) xor d(820) xor d(819) xor d(814) xor d(813) xor d(811) xor d(810) xor d(809) xor d(808) xor d(807) xor d(806) xor d(805) xor d(804) xor d(803) xor d(802) xor d(801) xor d(799) xor d(798) xor d(797) xor d(795) xor d(793) xor d(788) xor d(786) xor d(783) xor d(781) xor d(780) xor d(779) xor d(777) xor d(775) xor d(771) xor d(769) xor d(764) xor d(762) xor d(760) xor d(758) xor d(757) xor d(753) xor d(751) xor d(750) xor d(748) xor d(745) xor d(743) xor d(742) xor d(739) xor d(737) xor d(736) xor d(735) xor d(731) xor d(727) xor d(726) xor d(724) xor d(722) xor d(720) xor d(719) xor d(718) xor d(717) xor d(716) xor d(715) xor d(714) xor d(710) xor d(705) xor d(703) xor d(702) xor d(699) xor d(697) xor d(696) xor d(695) xor d(693) xor d(690) xor d(689) xor d(688) xor d(686) xor d(684) xor d(682) xor d(681) xor d(675) xor d(670) xor d(669) xor d(668) xor d(667) xor d(665) xor d(664) xor d(663) xor d(662) xor d(661) xor d(660) xor d(653) xor d(651) xor d(650) xor d(648) xor d(647) xor d(644) xor d(643) xor d(641) xor d(639) xor d(637) xor d(635) xor d(631) xor d(627) xor d(625) xor d(624) xor d(621) xor d(619) xor d(618) xor d(615) xor d(614) xor d(612) xor d(610) xor d(608) xor d(607) xor d(606) xor d(605) xor d(604) xor d(602) xor d(601) xor d(599) xor d(598) xor d(597) xor d(595) xor d(594) xor d(591) xor d(590) xor d(588) xor d(587) xor d(586) xor d(582) xor d(581) xor d(580) xor d(578) xor d(575) xor d(573) xor d(570) xor d(569) xor d(568) xor d(566) xor d(562) xor d(560) xor d(558) xor d(556) xor d(555) xor d(553) xor d(552) xor d(551) xor d(550) xor d(549) xor d(546) xor d(544) xor d(540) xor d(537) xor d(535) xor d(534) xor d(530) xor d(529) xor d(527) xor d(526) xor d(525) xor d(524) xor d(523) xor d(521) xor d(520) xor d(517) xor d(516) xor d(514) xor d(513) xor d(511) xor d(509) xor d(507) xor d(506) xor d(505) xor d(503) xor d(502) xor d(501) xor d(497) xor d(496) xor d(495) xor d(490) xor d(489) xor d(488) xor d(487) xor d(486) xor d(485) xor d(484) xor d(483) xor d(481) xor d(478) xor d(477) xor d(476) xor d(475) xor d(474) xor d(472) xor d(471) xor d(467) xor d(465) xor d(463) xor d(460) xor d(459) xor d(457) xor d(456) xor d(453) xor d(447) xor d(445) xor d(444) xor d(443) xor d(439) xor d(432) xor d(431) xor d(429) xor d(428) xor d(419) xor d(417) xor d(414) xor d(413) xor d(411) xor d(409) xor d(407) xor d(404) xor d(403) xor d(402) xor d(400) xor d(399) xor d(395) xor d(394) xor d(393) xor d(391) xor d(388) xor d(387) xor d(386) xor d(385) xor d(383) xor d(382) xor d(381) xor d(376) xor d(373) xor d(371) xor d(369) xor d(367) xor d(364) xor d(363) xor d(361) xor d(358) xor d(357) xor d(354) xor d(353) xor d(352) xor d(348) xor d(344) xor d(343) xor d(342) xor d(340) xor d(339) xor d(337) xor d(336) xor d(334) xor d(333) xor d(332) xor d(330) xor d(329) xor d(328) xor d(323) xor d(322) xor d(317) xor d(316) xor d(315) xor d(314) xor d(313) xor d(312) xor d(310) xor d(307) xor d(305) xor d(304) xor d(300) xor d(298) xor d(297) xor d(295) xor d(294) xor d(293) xor d(292) xor d(291) xor d(290) xor d(289) xor d(287) xor d(285) xor d(283) xor d(282) xor d(281) xor d(278) xor d(274) xor d(272) xor d(271) xor d(269) xor d(268) xor d(264) xor d(263) xor d(260) xor d(259) xor d(256) xor d(254) xor d(252) xor d(250) xor d(247) xor d(243) xor d(238) xor d(232) xor d(229) xor d(225) xor d(223) xor d(222) xor d(221) xor d(219) xor d(211) xor d(209) xor d(207) xor d(205) xor d(204) xor d(203) xor d(202) xor d(198) xor d(197) xor d(196) xor d(194) xor d(193) xor d(192) xor d(189) xor d(188) xor d(187) xor d(186) xor d(185) xor d(183) xor d(181) xor d(178) xor d(177) xor d(167) xor d(166) xor d(165) xor d(164) xor d(162) xor d(161) xor d(157) xor d(156) xor d(153) xor d(151) xor d(150) xor d(146) xor d(144) xor d(139) xor d(138) xor d(132) xor d(131) xor d(130) xor d(129) xor d(127) xor d(123) xor d(122) xor d(121) xor d(120) xor d(118) xor d(114) xor d(113) xor d(112) xor d(111) xor d(109) xor d(108) xor d(106) xor d(105) xor d(101) xor d(99) xor d(98) xor d(96) xor d(94) xor d(93) xor d(92) xor d(91) xor d(90) xor d(89) xor d(82) xor d(80) xor d(79) xor d(78) xor d(77) xor d(76) xor d(74) xor d(68) xor d(67) xor d(63) xor d(62) xor d(61) xor d(60) xor d(58) xor d(56) xor d(55) xor d(53) xor d(50) xor d(49) xor d(48) xor d(45) xor d(43) xor d(42) xor d(40) xor d(39) xor d(32) xor d(29) xor d(27) xor d(26) xor d(25) xor d(24) xor d(23) xor d(21) xor d(20) xor d(19) xor d(11) xor d(7) xor d(5) xor d(4) xor d(1) xor c(1) xor c(2) xor c(3) xor c(7) xor c(8) xor c(9) xor c(11) xor c(12) xor c(14) xor c(15) xor c(18) xor c(19) xor c(21) xor c(22) xor c(24) xor c(27) xor c(28) xor c(31);
    newcrc(28) := d(1021) xor d(1020) xor d(1017) xor d(1015) xor d(1014) xor d(1012) xor d(1011) xor d(1008) xor d(1007) xor d(1005) xor d(1004) xor d(1002) xor d(1001) xor d(1000) xor d(996) xor d(995) xor d(994) xor d(992) xor d(990) xor d(988) xor d(986) xor d(981) xor d(980) xor d(979) xor d(978) xor d(977) xor d(976) xor d(975) xor d(974) xor d(973) xor d(971) xor d(970) xor d(967) xor d(963) xor d(956) xor d(955) xor d(954) xor d(951) xor d(950) xor d(949) xor d(946) xor d(944) xor d(940) xor d(937) xor d(935) xor d(934) xor d(931) xor d(930) xor d(929) xor d(927) xor d(916) xor d(914) xor d(913) xor d(911) xor d(906) xor d(903) xor d(902) xor d(900) xor d(899) xor d(898) xor d(897) xor d(896) xor d(895) xor d(894) xor d(893) xor d(892) xor d(889) xor d(887) xor d(886) xor d(885) xor d(883) xor d(882) xor d(879) xor d(877) xor d(875) xor d(874) xor d(873) xor d(872) xor d(871) xor d(870) xor d(869) xor d(867) xor d(865) xor d(864) xor d(863) xor d(859) xor d(857) xor d(856) xor d(855) xor d(853) xor d(850) xor d(849) xor d(847) xor d(846) xor d(845) xor d(844) xor d(842) xor d(838) xor d(836) xor d(835) xor d(833) xor d(831) xor d(830) xor d(828) xor d(823) xor d(821) xor d(820) xor d(815) xor d(814) xor d(812) xor d(811) xor d(810) xor d(809) xor d(808) xor d(807) xor d(806) xor d(805) xor d(804) xor d(803) xor d(802) xor d(800) xor d(799) xor d(798) xor d(796) xor d(794) xor d(789) xor d(787) xor d(784) xor d(782) xor d(781) xor d(780) xor d(778) xor d(776) xor d(772) xor d(770) xor d(765) xor d(763) xor d(761) xor d(759) xor d(758) xor d(754) xor d(752) xor d(751) xor d(749) xor d(746) xor d(744) xor d(743) xor d(740) xor d(738) xor d(737) xor d(736) xor d(732) xor d(728) xor d(727) xor d(725) xor d(723) xor d(721) xor d(720) xor d(719) xor d(718) xor d(717) xor d(716) xor d(715) xor d(711) xor d(706) xor d(704) xor d(703) xor d(700) xor d(698) xor d(697) xor d(696) xor d(694) xor d(691) xor d(690) xor d(689) xor d(687) xor d(685) xor d(683) xor d(682) xor d(676) xor d(671) xor d(670) xor d(669) xor d(668) xor d(666) xor d(665) xor d(664) xor d(663) xor d(662) xor d(661) xor d(654) xor d(652) xor d(651) xor d(649) xor d(648) xor d(645) xor d(644) xor d(642) xor d(640) xor d(638) xor d(636) xor d(632) xor d(628) xor d(626) xor d(625) xor d(622) xor d(620) xor d(619) xor d(616) xor d(615) xor d(613) xor d(611) xor d(609) xor d(608) xor d(607) xor d(606) xor d(605) xor d(603) xor d(602) xor d(600) xor d(599) xor d(598) xor d(596) xor d(595) xor d(592) xor d(591) xor d(589) xor d(588) xor d(587) xor d(583) xor d(582) xor d(581) xor d(579) xor d(576) xor d(574) xor d(571) xor d(570) xor d(569) xor d(567) xor d(563) xor d(561) xor d(559) xor d(557) xor d(556) xor d(554) xor d(553) xor d(552) xor d(551) xor d(550) xor d(547) xor d(545) xor d(541) xor d(538) xor d(536) xor d(535) xor d(531) xor d(530) xor d(528) xor d(527) xor d(526) xor d(525) xor d(524) xor d(522) xor d(521) xor d(518) xor d(517) xor d(515) xor d(514) xor d(512) xor d(510) xor d(508) xor d(507) xor d(506) xor d(504) xor d(503) xor d(502) xor d(498) xor d(497) xor d(496) xor d(491) xor d(490) xor d(489) xor d(488) xor d(487) xor d(486) xor d(485) xor d(484) xor d(482) xor d(479) xor d(478) xor d(477) xor d(476) xor d(475) xor d(473) xor d(472) xor d(468) xor d(466) xor d(464) xor d(461) xor d(460) xor d(458) xor d(457) xor d(454) xor d(448) xor d(446) xor d(445) xor d(444) xor d(440) xor d(433) xor d(432) xor d(430) xor d(429) xor d(420) xor d(418) xor d(415) xor d(414) xor d(412) xor d(410) xor d(408) xor d(405) xor d(404) xor d(403) xor d(401) xor d(400) xor d(396) xor d(395) xor d(394) xor d(392) xor d(389) xor d(388) xor d(387) xor d(386) xor d(384) xor d(383) xor d(382) xor d(377) xor d(374) xor d(372) xor d(370) xor d(368) xor d(365) xor d(364) xor d(362) xor d(359) xor d(358) xor d(355) xor d(354) xor d(353) xor d(349) xor d(345) xor d(344) xor d(343) xor d(341) xor d(340) xor d(338) xor d(337) xor d(335) xor d(334) xor d(333) xor d(331) xor d(330) xor d(329) xor d(324) xor d(323) xor d(318) xor d(317) xor d(316) xor d(315) xor d(314) xor d(313) xor d(311) xor d(308) xor d(306) xor d(305) xor d(301) xor d(299) xor d(298) xor d(296) xor d(295) xor d(294) xor d(293) xor d(292) xor d(291) xor d(290) xor d(288) xor d(286) xor d(284) xor d(283) xor d(282) xor d(279) xor d(275) xor d(273) xor d(272) xor d(270) xor d(269) xor d(265) xor d(264) xor d(261) xor d(260) xor d(257) xor d(255) xor d(253) xor d(251) xor d(248) xor d(244) xor d(239) xor d(233) xor d(230) xor d(226) xor d(224) xor d(223) xor d(222) xor d(220) xor d(212) xor d(210) xor d(208) xor d(206) xor d(205) xor d(204) xor d(203) xor d(199) xor d(198) xor d(197) xor d(195) xor d(194) xor d(193) xor d(190) xor d(189) xor d(188) xor d(187) xor d(186) xor d(184) xor d(182) xor d(179) xor d(178) xor d(168) xor d(167) xor d(166) xor d(165) xor d(163) xor d(162) xor d(158) xor d(157) xor d(154) xor d(152) xor d(151) xor d(147) xor d(145) xor d(140) xor d(139) xor d(133) xor d(132) xor d(131) xor d(130) xor d(128) xor d(124) xor d(123) xor d(122) xor d(121) xor d(119) xor d(115) xor d(114) xor d(113) xor d(112) xor d(110) xor d(109) xor d(107) xor d(106) xor d(102) xor d(100) xor d(99) xor d(97) xor d(95) xor d(94) xor d(93) xor d(92) xor d(91) xor d(90) xor d(83) xor d(81) xor d(80) xor d(79) xor d(78) xor d(77) xor d(75) xor d(69) xor d(68) xor d(64) xor d(63) xor d(62) xor d(61) xor d(59) xor d(57) xor d(56) xor d(54) xor d(51) xor d(50) xor d(49) xor d(46) xor d(44) xor d(43) xor d(41) xor d(40) xor d(33) xor d(30) xor d(28) xor d(27) xor d(26) xor d(25) xor d(24) xor d(22) xor d(21) xor d(20) xor d(12) xor d(8) xor d(6) xor d(5) xor d(2) xor c(0) xor c(2) xor c(3) xor c(4) xor c(8) xor c(9) xor c(10) xor c(12) xor c(13) xor c(15) xor c(16) xor c(19) xor c(20) xor c(22) xor c(23) xor c(25) xor c(28) xor c(29);
    newcrc(29) := d(1022) xor d(1021) xor d(1018) xor d(1016) xor d(1015) xor d(1013) xor d(1012) xor d(1009) xor d(1008) xor d(1006) xor d(1005) xor d(1003) xor d(1002) xor d(1001) xor d(997) xor d(996) xor d(995) xor d(993) xor d(991) xor d(989) xor d(987) xor d(982) xor d(981) xor d(980) xor d(979) xor d(978) xor d(977) xor d(976) xor d(975) xor d(974) xor d(972) xor d(971) xor d(968) xor d(964) xor d(957) xor d(956) xor d(955) xor d(952) xor d(951) xor d(950) xor d(947) xor d(945) xor d(941) xor d(938) xor d(936) xor d(935) xor d(932) xor d(931) xor d(930) xor d(928) xor d(917) xor d(915) xor d(914) xor d(912) xor d(907) xor d(904) xor d(903) xor d(901) xor d(900) xor d(899) xor d(898) xor d(897) xor d(896) xor d(895) xor d(894) xor d(893) xor d(890) xor d(888) xor d(887) xor d(886) xor d(884) xor d(883) xor d(880) xor d(878) xor d(876) xor d(875) xor d(874) xor d(873) xor d(872) xor d(871) xor d(870) xor d(868) xor d(866) xor d(865) xor d(864) xor d(860) xor d(858) xor d(857) xor d(856) xor d(854) xor d(851) xor d(850) xor d(848) xor d(847) xor d(846) xor d(845) xor d(843) xor d(839) xor d(837) xor d(836) xor d(834) xor d(832) xor d(831) xor d(829) xor d(824) xor d(822) xor d(821) xor d(816) xor d(815) xor d(813) xor d(812) xor d(811) xor d(810) xor d(809) xor d(808) xor d(807) xor d(806) xor d(805) xor d(804) xor d(803) xor d(801) xor d(800) xor d(799) xor d(797) xor d(795) xor d(790) xor d(788) xor d(785) xor d(783) xor d(782) xor d(781) xor d(779) xor d(777) xor d(773) xor d(771) xor d(766) xor d(764) xor d(762) xor d(760) xor d(759) xor d(755) xor d(753) xor d(752) xor d(750) xor d(747) xor d(745) xor d(744) xor d(741) xor d(739) xor d(738) xor d(737) xor d(733) xor d(729) xor d(728) xor d(726) xor d(724) xor d(722) xor d(721) xor d(720) xor d(719) xor d(718) xor d(717) xor d(716) xor d(712) xor d(707) xor d(705) xor d(704) xor d(701) xor d(699) xor d(698) xor d(697) xor d(695) xor d(692) xor d(691) xor d(690) xor d(688) xor d(686) xor d(684) xor d(683) xor d(677) xor d(672) xor d(671) xor d(670) xor d(669) xor d(667) xor d(666) xor d(665) xor d(664) xor d(663) xor d(662) xor d(655) xor d(653) xor d(652) xor d(650) xor d(649) xor d(646) xor d(645) xor d(643) xor d(641) xor d(639) xor d(637) xor d(633) xor d(629) xor d(627) xor d(626) xor d(623) xor d(621) xor d(620) xor d(617) xor d(616) xor d(614) xor d(612) xor d(610) xor d(609) xor d(608) xor d(607) xor d(606) xor d(604) xor d(603) xor d(601) xor d(600) xor d(599) xor d(597) xor d(596) xor d(593) xor d(592) xor d(590) xor d(589) xor d(588) xor d(584) xor d(583) xor d(582) xor d(580) xor d(577) xor d(575) xor d(572) xor d(571) xor d(570) xor d(568) xor d(564) xor d(562) xor d(560) xor d(558) xor d(557) xor d(555) xor d(554) xor d(553) xor d(552) xor d(551) xor d(548) xor d(546) xor d(542) xor d(539) xor d(537) xor d(536) xor d(532) xor d(531) xor d(529) xor d(528) xor d(527) xor d(526) xor d(525) xor d(523) xor d(522) xor d(519) xor d(518) xor d(516) xor d(515) xor d(513) xor d(511) xor d(509) xor d(508) xor d(507) xor d(505) xor d(504) xor d(503) xor d(499) xor d(498) xor d(497) xor d(492) xor d(491) xor d(490) xor d(489) xor d(488) xor d(487) xor d(486) xor d(485) xor d(483) xor d(480) xor d(479) xor d(478) xor d(477) xor d(476) xor d(474) xor d(473) xor d(469) xor d(467) xor d(465) xor d(462) xor d(461) xor d(459) xor d(458) xor d(455) xor d(449) xor d(447) xor d(446) xor d(445) xor d(441) xor d(434) xor d(433) xor d(431) xor d(430) xor d(421) xor d(419) xor d(416) xor d(415) xor d(413) xor d(411) xor d(409) xor d(406) xor d(405) xor d(404) xor d(402) xor d(401) xor d(397) xor d(396) xor d(395) xor d(393) xor d(390) xor d(389) xor d(388) xor d(387) xor d(385) xor d(384) xor d(383) xor d(378) xor d(375) xor d(373) xor d(371) xor d(369) xor d(366) xor d(365) xor d(363) xor d(360) xor d(359) xor d(356) xor d(355) xor d(354) xor d(350) xor d(346) xor d(345) xor d(344) xor d(342) xor d(341) xor d(339) xor d(338) xor d(336) xor d(335) xor d(334) xor d(332) xor d(331) xor d(330) xor d(325) xor d(324) xor d(319) xor d(318) xor d(317) xor d(316) xor d(315) xor d(314) xor d(312) xor d(309) xor d(307) xor d(306) xor d(302) xor d(300) xor d(299) xor d(297) xor d(296) xor d(295) xor d(294) xor d(293) xor d(292) xor d(291) xor d(289) xor d(287) xor d(285) xor d(284) xor d(283) xor d(280) xor d(276) xor d(274) xor d(273) xor d(271) xor d(270) xor d(266) xor d(265) xor d(262) xor d(261) xor d(258) xor d(256) xor d(254) xor d(252) xor d(249) xor d(245) xor d(240) xor d(234) xor d(231) xor d(227) xor d(225) xor d(224) xor d(223) xor d(221) xor d(213) xor d(211) xor d(209) xor d(207) xor d(206) xor d(205) xor d(204) xor d(200) xor d(199) xor d(198) xor d(196) xor d(195) xor d(194) xor d(191) xor d(190) xor d(189) xor d(188) xor d(187) xor d(185) xor d(183) xor d(180) xor d(179) xor d(169) xor d(168) xor d(167) xor d(166) xor d(164) xor d(163) xor d(159) xor d(158) xor d(155) xor d(153) xor d(152) xor d(148) xor d(146) xor d(141) xor d(140) xor d(134) xor d(133) xor d(132) xor d(131) xor d(129) xor d(125) xor d(124) xor d(123) xor d(122) xor d(120) xor d(116) xor d(115) xor d(114) xor d(113) xor d(111) xor d(110) xor d(108) xor d(107) xor d(103) xor d(101) xor d(100) xor d(98) xor d(96) xor d(95) xor d(94) xor d(93) xor d(92) xor d(91) xor d(84) xor d(82) xor d(81) xor d(80) xor d(79) xor d(78) xor d(76) xor d(70) xor d(69) xor d(65) xor d(64) xor d(63) xor d(62) xor d(60) xor d(58) xor d(57) xor d(55) xor d(52) xor d(51) xor d(50) xor d(47) xor d(45) xor d(44) xor d(42) xor d(41) xor d(34) xor d(31) xor d(29) xor d(28) xor d(27) xor d(26) xor d(25) xor d(23) xor d(22) xor d(21) xor d(13) xor d(9) xor d(7) xor d(6) xor d(3) xor c(1) xor c(3) xor c(4) xor c(5) xor c(9) xor c(10) xor c(11) xor c(13) xor c(14) xor c(16) xor c(17) xor c(20) xor c(21) xor c(23) xor c(24) xor c(26) xor c(29) xor c(30);
    newcrc(30) := d(1023) xor d(1022) xor d(1019) xor d(1017) xor d(1016) xor d(1014) xor d(1013) xor d(1010) xor d(1009) xor d(1007) xor d(1006) xor d(1004) xor d(1003) xor d(1002) xor d(998) xor d(997) xor d(996) xor d(994) xor d(992) xor d(990) xor d(988) xor d(983) xor d(982) xor d(981) xor d(980) xor d(979) xor d(978) xor d(977) xor d(976) xor d(975) xor d(973) xor d(972) xor d(969) xor d(965) xor d(958) xor d(957) xor d(956) xor d(953) xor d(952) xor d(951) xor d(948) xor d(946) xor d(942) xor d(939) xor d(937) xor d(936) xor d(933) xor d(932) xor d(931) xor d(929) xor d(918) xor d(916) xor d(915) xor d(913) xor d(908) xor d(905) xor d(904) xor d(902) xor d(901) xor d(900) xor d(899) xor d(898) xor d(897) xor d(896) xor d(895) xor d(894) xor d(891) xor d(889) xor d(888) xor d(887) xor d(885) xor d(884) xor d(881) xor d(879) xor d(877) xor d(876) xor d(875) xor d(874) xor d(873) xor d(872) xor d(871) xor d(869) xor d(867) xor d(866) xor d(865) xor d(861) xor d(859) xor d(858) xor d(857) xor d(855) xor d(852) xor d(851) xor d(849) xor d(848) xor d(847) xor d(846) xor d(844) xor d(840) xor d(838) xor d(837) xor d(835) xor d(833) xor d(832) xor d(830) xor d(825) xor d(823) xor d(822) xor d(817) xor d(816) xor d(814) xor d(813) xor d(812) xor d(811) xor d(810) xor d(809) xor d(808) xor d(807) xor d(806) xor d(805) xor d(804) xor d(802) xor d(801) xor d(800) xor d(798) xor d(796) xor d(791) xor d(789) xor d(786) xor d(784) xor d(783) xor d(782) xor d(780) xor d(778) xor d(774) xor d(772) xor d(767) xor d(765) xor d(763) xor d(761) xor d(760) xor d(756) xor d(754) xor d(753) xor d(751) xor d(748) xor d(746) xor d(745) xor d(742) xor d(740) xor d(739) xor d(738) xor d(734) xor d(730) xor d(729) xor d(727) xor d(725) xor d(723) xor d(722) xor d(721) xor d(720) xor d(719) xor d(718) xor d(717) xor d(713) xor d(708) xor d(706) xor d(705) xor d(702) xor d(700) xor d(699) xor d(698) xor d(696) xor d(693) xor d(692) xor d(691) xor d(689) xor d(687) xor d(685) xor d(684) xor d(678) xor d(673) xor d(672) xor d(671) xor d(670) xor d(668) xor d(667) xor d(666) xor d(665) xor d(664) xor d(663) xor d(656) xor d(654) xor d(653) xor d(651) xor d(650) xor d(647) xor d(646) xor d(644) xor d(642) xor d(640) xor d(638) xor d(634) xor d(630) xor d(628) xor d(627) xor d(624) xor d(622) xor d(621) xor d(618) xor d(617) xor d(615) xor d(613) xor d(611) xor d(610) xor d(609) xor d(608) xor d(607) xor d(605) xor d(604) xor d(602) xor d(601) xor d(600) xor d(598) xor d(597) xor d(594) xor d(593) xor d(591) xor d(590) xor d(589) xor d(585) xor d(584) xor d(583) xor d(581) xor d(578) xor d(576) xor d(573) xor d(572) xor d(571) xor d(569) xor d(565) xor d(563) xor d(561) xor d(559) xor d(558) xor d(556) xor d(555) xor d(554) xor d(553) xor d(552) xor d(549) xor d(547) xor d(543) xor d(540) xor d(538) xor d(537) xor d(533) xor d(532) xor d(530) xor d(529) xor d(528) xor d(527) xor d(526) xor d(524) xor d(523) xor d(520) xor d(519) xor d(517) xor d(516) xor d(514) xor d(512) xor d(510) xor d(509) xor d(508) xor d(506) xor d(505) xor d(504) xor d(500) xor d(499) xor d(498) xor d(493) xor d(492) xor d(491) xor d(490) xor d(489) xor d(488) xor d(487) xor d(486) xor d(484) xor d(481) xor d(480) xor d(479) xor d(478) xor d(477) xor d(475) xor d(474) xor d(470) xor d(468) xor d(466) xor d(463) xor d(462) xor d(460) xor d(459) xor d(456) xor d(450) xor d(448) xor d(447) xor d(446) xor d(442) xor d(435) xor d(434) xor d(432) xor d(431) xor d(422) xor d(420) xor d(417) xor d(416) xor d(414) xor d(412) xor d(410) xor d(407) xor d(406) xor d(405) xor d(403) xor d(402) xor d(398) xor d(397) xor d(396) xor d(394) xor d(391) xor d(390) xor d(389) xor d(388) xor d(386) xor d(385) xor d(384) xor d(379) xor d(376) xor d(374) xor d(372) xor d(370) xor d(367) xor d(366) xor d(364) xor d(361) xor d(360) xor d(357) xor d(356) xor d(355) xor d(351) xor d(347) xor d(346) xor d(345) xor d(343) xor d(342) xor d(340) xor d(339) xor d(337) xor d(336) xor d(335) xor d(333) xor d(332) xor d(331) xor d(326) xor d(325) xor d(320) xor d(319) xor d(318) xor d(317) xor d(316) xor d(315) xor d(313) xor d(310) xor d(308) xor d(307) xor d(303) xor d(301) xor d(300) xor d(298) xor d(297) xor d(296) xor d(295) xor d(294) xor d(293) xor d(292) xor d(290) xor d(288) xor d(286) xor d(285) xor d(284) xor d(281) xor d(277) xor d(275) xor d(274) xor d(272) xor d(271) xor d(267) xor d(266) xor d(263) xor d(262) xor d(259) xor d(257) xor d(255) xor d(253) xor d(250) xor d(246) xor d(241) xor d(235) xor d(232) xor d(228) xor d(226) xor d(225) xor d(224) xor d(222) xor d(214) xor d(212) xor d(210) xor d(208) xor d(207) xor d(206) xor d(205) xor d(201) xor d(200) xor d(199) xor d(197) xor d(196) xor d(195) xor d(192) xor d(191) xor d(190) xor d(189) xor d(188) xor d(186) xor d(184) xor d(181) xor d(180) xor d(170) xor d(169) xor d(168) xor d(167) xor d(165) xor d(164) xor d(160) xor d(159) xor d(156) xor d(154) xor d(153) xor d(149) xor d(147) xor d(142) xor d(141) xor d(135) xor d(134) xor d(133) xor d(132) xor d(130) xor d(126) xor d(125) xor d(124) xor d(123) xor d(121) xor d(117) xor d(116) xor d(115) xor d(114) xor d(112) xor d(111) xor d(109) xor d(108) xor d(104) xor d(102) xor d(101) xor d(99) xor d(97) xor d(96) xor d(95) xor d(94) xor d(93) xor d(92) xor d(85) xor d(83) xor d(82) xor d(81) xor d(80) xor d(79) xor d(77) xor d(71) xor d(70) xor d(66) xor d(65) xor d(64) xor d(63) xor d(61) xor d(59) xor d(58) xor d(56) xor d(53) xor d(52) xor d(51) xor d(48) xor d(46) xor d(45) xor d(43) xor d(42) xor d(35) xor d(32) xor d(30) xor d(29) xor d(28) xor d(27) xor d(26) xor d(24) xor d(23) xor d(22) xor d(14) xor d(10) xor d(8) xor d(7) xor d(4) xor c(0) xor c(2) xor c(4) xor c(5) xor c(6) xor c(10) xor c(11) xor c(12) xor c(14) xor c(15) xor c(17) xor c(18) xor c(21) xor c(22) xor c(24) xor c(25) xor c(27) xor c(30) xor c(31);
    newcrc(31) := d(1023) xor d(1020) xor d(1018) xor d(1017) xor d(1015) xor d(1014) xor d(1011) xor d(1010) xor d(1008) xor d(1007) xor d(1005) xor d(1004) xor d(1003) xor d(999) xor d(998) xor d(997) xor d(995) xor d(993) xor d(991) xor d(989) xor d(984) xor d(983) xor d(982) xor d(981) xor d(980) xor d(979) xor d(978) xor d(977) xor d(976) xor d(974) xor d(973) xor d(970) xor d(966) xor d(959) xor d(958) xor d(957) xor d(954) xor d(953) xor d(952) xor d(949) xor d(947) xor d(943) xor d(940) xor d(938) xor d(937) xor d(934) xor d(933) xor d(932) xor d(930) xor d(919) xor d(917) xor d(916) xor d(914) xor d(909) xor d(906) xor d(905) xor d(903) xor d(902) xor d(901) xor d(900) xor d(899) xor d(898) xor d(897) xor d(896) xor d(895) xor d(892) xor d(890) xor d(889) xor d(888) xor d(886) xor d(885) xor d(882) xor d(880) xor d(878) xor d(877) xor d(876) xor d(875) xor d(874) xor d(873) xor d(872) xor d(870) xor d(868) xor d(867) xor d(866) xor d(862) xor d(860) xor d(859) xor d(858) xor d(856) xor d(853) xor d(852) xor d(850) xor d(849) xor d(848) xor d(847) xor d(845) xor d(841) xor d(839) xor d(838) xor d(836) xor d(834) xor d(833) xor d(831) xor d(826) xor d(824) xor d(823) xor d(818) xor d(817) xor d(815) xor d(814) xor d(813) xor d(812) xor d(811) xor d(810) xor d(809) xor d(808) xor d(807) xor d(806) xor d(805) xor d(803) xor d(802) xor d(801) xor d(799) xor d(797) xor d(792) xor d(790) xor d(787) xor d(785) xor d(784) xor d(783) xor d(781) xor d(779) xor d(775) xor d(773) xor d(768) xor d(766) xor d(764) xor d(762) xor d(761) xor d(757) xor d(755) xor d(754) xor d(752) xor d(749) xor d(747) xor d(746) xor d(743) xor d(741) xor d(740) xor d(739) xor d(735) xor d(731) xor d(730) xor d(728) xor d(726) xor d(724) xor d(723) xor d(722) xor d(721) xor d(720) xor d(719) xor d(718) xor d(714) xor d(709) xor d(707) xor d(706) xor d(703) xor d(701) xor d(700) xor d(699) xor d(697) xor d(694) xor d(693) xor d(692) xor d(690) xor d(688) xor d(686) xor d(685) xor d(679) xor d(674) xor d(673) xor d(672) xor d(671) xor d(669) xor d(668) xor d(667) xor d(666) xor d(665) xor d(664) xor d(657) xor d(655) xor d(654) xor d(652) xor d(651) xor d(648) xor d(647) xor d(645) xor d(643) xor d(641) xor d(639) xor d(635) xor d(631) xor d(629) xor d(628) xor d(625) xor d(623) xor d(622) xor d(619) xor d(618) xor d(616) xor d(614) xor d(612) xor d(611) xor d(610) xor d(609) xor d(608) xor d(606) xor d(605) xor d(603) xor d(602) xor d(601) xor d(599) xor d(598) xor d(595) xor d(594) xor d(592) xor d(591) xor d(590) xor d(586) xor d(585) xor d(584) xor d(582) xor d(579) xor d(577) xor d(574) xor d(573) xor d(572) xor d(570) xor d(566) xor d(564) xor d(562) xor d(560) xor d(559) xor d(557) xor d(556) xor d(555) xor d(554) xor d(553) xor d(550) xor d(548) xor d(544) xor d(541) xor d(539) xor d(538) xor d(534) xor d(533) xor d(531) xor d(530) xor d(529) xor d(528) xor d(527) xor d(525) xor d(524) xor d(521) xor d(520) xor d(518) xor d(517) xor d(515) xor d(513) xor d(511) xor d(510) xor d(509) xor d(507) xor d(506) xor d(505) xor d(501) xor d(500) xor d(499) xor d(494) xor d(493) xor d(492) xor d(491) xor d(490) xor d(489) xor d(488) xor d(487) xor d(485) xor d(482) xor d(481) xor d(480) xor d(479) xor d(478) xor d(476) xor d(475) xor d(471) xor d(469) xor d(467) xor d(464) xor d(463) xor d(461) xor d(460) xor d(457) xor d(451) xor d(449) xor d(448) xor d(447) xor d(443) xor d(436) xor d(435) xor d(433) xor d(432) xor d(423) xor d(421) xor d(418) xor d(417) xor d(415) xor d(413) xor d(411) xor d(408) xor d(407) xor d(406) xor d(404) xor d(403) xor d(399) xor d(398) xor d(397) xor d(395) xor d(392) xor d(391) xor d(390) xor d(389) xor d(387) xor d(386) xor d(385) xor d(380) xor d(377) xor d(375) xor d(373) xor d(371) xor d(368) xor d(367) xor d(365) xor d(362) xor d(361) xor d(358) xor d(357) xor d(356) xor d(352) xor d(348) xor d(347) xor d(346) xor d(344) xor d(343) xor d(341) xor d(340) xor d(338) xor d(337) xor d(336) xor d(334) xor d(333) xor d(332) xor d(327) xor d(326) xor d(321) xor d(320) xor d(319) xor d(318) xor d(317) xor d(316) xor d(314) xor d(311) xor d(309) xor d(308) xor d(304) xor d(302) xor d(301) xor d(299) xor d(298) xor d(297) xor d(296) xor d(295) xor d(294) xor d(293) xor d(291) xor d(289) xor d(287) xor d(286) xor d(285) xor d(282) xor d(278) xor d(276) xor d(275) xor d(273) xor d(272) xor d(268) xor d(267) xor d(264) xor d(263) xor d(260) xor d(258) xor d(256) xor d(254) xor d(251) xor d(247) xor d(242) xor d(236) xor d(233) xor d(229) xor d(227) xor d(226) xor d(225) xor d(223) xor d(215) xor d(213) xor d(211) xor d(209) xor d(208) xor d(207) xor d(206) xor d(202) xor d(201) xor d(200) xor d(198) xor d(197) xor d(196) xor d(193) xor d(192) xor d(191) xor d(190) xor d(189) xor d(187) xor d(185) xor d(182) xor d(181) xor d(171) xor d(170) xor d(169) xor d(168) xor d(166) xor d(165) xor d(161) xor d(160) xor d(157) xor d(155) xor d(154) xor d(150) xor d(148) xor d(143) xor d(142) xor d(136) xor d(135) xor d(134) xor d(133) xor d(131) xor d(127) xor d(126) xor d(125) xor d(124) xor d(122) xor d(118) xor d(117) xor d(116) xor d(115) xor d(113) xor d(112) xor d(110) xor d(109) xor d(105) xor d(103) xor d(102) xor d(100) xor d(98) xor d(97) xor d(96) xor d(95) xor d(94) xor d(93) xor d(86) xor d(84) xor d(83) xor d(82) xor d(81) xor d(80) xor d(78) xor d(72) xor d(71) xor d(67) xor d(66) xor d(65) xor d(64) xor d(62) xor d(60) xor d(59) xor d(57) xor d(54) xor d(53) xor d(52) xor d(49) xor d(47) xor d(46) xor d(44) xor d(43) xor d(36) xor d(33) xor d(31) xor d(30) xor d(29) xor d(28) xor d(27) xor d(25) xor d(24) xor d(23) xor d(15) xor d(11) xor d(9) xor d(8) xor d(5) xor c(1) xor c(3) xor c(5) xor c(6) xor c(7) xor c(11) xor c(12) xor c(13) xor c(15) xor c(16) xor c(18) xor c(19) xor c(22) xor c(23) xor c(25) xor c(26) xor c(28) xor c(31);
    return newcrc;
  end nextCRC32_D1024;

end PCK_CRC32_D1024;
